--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.10.03 (64-bit)
--Part Number: GW2A-LV18PG256C8/I7
--Device: GW2A-18
--Device Version: C
--Created Time: Mon Nov 18 12:53:53 2024

library IEEE;
use IEEE.std_logic_1164.all;

entity vga_sample_buf is
    port (
        douta: out std_logic_vector(17 downto 0);
        doutb: out std_logic_vector(17 downto 0);
        clka: in std_logic;
        ocea: in std_logic;
        cea: in std_logic;
        reseta: in std_logic;
        wrea: in std_logic;
        clkb: in std_logic;
        oceb: in std_logic;
        ceb: in std_logic;
        resetb: in std_logic;
        wreb: in std_logic;
        ada: in std_logic_vector(10 downto 0);
        dina: in std_logic_vector(17 downto 0);
        adb: in std_logic_vector(10 downto 0);
        dinb: in std_logic_vector(17 downto 0)
    );
end vga_sample_buf;

architecture Behavioral of vga_sample_buf is

    signal dpx9b_inst_0_douta_w: std_logic_vector(8 downto 0);
    signal dpx9b_inst_0_doutb_w: std_logic_vector(8 downto 0);
    signal dpx9b_inst_1_douta_w: std_logic_vector(8 downto 0);
    signal dpx9b_inst_1_doutb_w: std_logic_vector(8 downto 0);
    signal gw_gnd: std_logic;
    signal dpx9b_inst_0_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpx9b_inst_0_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpx9b_inst_0_ADA_i: std_logic_vector(13 downto 0);
    signal dpx9b_inst_0_DIA_i: std_logic_vector(17 downto 0);
    signal dpx9b_inst_0_ADB_i: std_logic_vector(13 downto 0);
    signal dpx9b_inst_0_DIB_i: std_logic_vector(17 downto 0);
    signal dpx9b_inst_0_DOA_o: std_logic_vector(17 downto 0);
    signal dpx9b_inst_0_DOB_o: std_logic_vector(17 downto 0);
    signal dpx9b_inst_1_BLKSELA_i: std_logic_vector(2 downto 0);
    signal dpx9b_inst_1_BLKSELB_i: std_logic_vector(2 downto 0);
    signal dpx9b_inst_1_ADA_i: std_logic_vector(13 downto 0);
    signal dpx9b_inst_1_DIA_i: std_logic_vector(17 downto 0);
    signal dpx9b_inst_1_ADB_i: std_logic_vector(13 downto 0);
    signal dpx9b_inst_1_DIB_i: std_logic_vector(17 downto 0);
    signal dpx9b_inst_1_DOA_o: std_logic_vector(17 downto 0);
    signal dpx9b_inst_1_DOB_o: std_logic_vector(17 downto 0);

    --component declaration
    component DPX9B
        generic (
            READ_MODE0: in bit := '0';
            READ_MODE1: in bit := '0';
            WRITE_MODE0: in bit_vector := "00";
            WRITE_MODE1: in bit_vector := "00";
            BIT_WIDTH_0: in integer :=18;
            BIT_WIDTH_1: in integer :=18;
            BLK_SEL_0: in bit_vector := "000";
            BLK_SEL_1: in bit_vector := "000";
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"000000000000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DOA: out std_logic_vector(17 downto 0);
            DOB: out std_logic_vector(17 downto 0);
            CLKA: in std_logic;
            OCEA: in std_logic;
            CEA: in std_logic;
            RESETA: in std_logic;
            WREA: in std_logic;
            CLKB: in std_logic;
            OCEB: in std_logic;
            CEB: in std_logic;
            RESETB: in std_logic;
            WREB: in std_logic;
            BLKSELA: in std_logic_vector(2 downto 0);
            BLKSELB: in std_logic_vector(2 downto 0);
            ADA: in std_logic_vector(13 downto 0);
            DIA: in std_logic_vector(17 downto 0);
            ADB: in std_logic_vector(13 downto 0);
            DIB: in std_logic_vector(17 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    dpx9b_inst_0_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_0_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_0_ADA_i <= ada(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_0_DIA_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & dina(8 downto 0);
    dpx9b_inst_0_ADB_i <= adb(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_0_DIB_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & dinb(8 downto 0);
    douta(8 downto 0) <= dpx9b_inst_0_DOA_o(8 downto 0) ;
    dpx9b_inst_0_douta_w(8 downto 0) <= dpx9b_inst_0_DOA_o(17 downto 9) ;
    doutb(8 downto 0) <= dpx9b_inst_0_DOB_o(8 downto 0) ;
    dpx9b_inst_0_doutb_w(8 downto 0) <= dpx9b_inst_0_DOB_o(17 downto 9) ;
    dpx9b_inst_1_BLKSELA_i <= gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_1_BLKSELB_i <= gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_1_ADA_i <= ada(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_1_DIA_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & dina(17 downto 9);
    dpx9b_inst_1_ADB_i <= adb(10 downto 0) & gw_gnd & gw_gnd & gw_gnd;
    dpx9b_inst_1_DIB_i <= gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & gw_gnd & dinb(17 downto 9);
    douta(17 downto 9) <= dpx9b_inst_1_DOA_o(8 downto 0) ;
    dpx9b_inst_1_douta_w(8 downto 0) <= dpx9b_inst_1_DOA_o(17 downto 9) ;
    doutb(17 downto 9) <= dpx9b_inst_1_DOB_o(8 downto 0) ;
    dpx9b_inst_1_doutb_w(8 downto 0) <= dpx9b_inst_1_DOB_o(17 downto 9) ;

    dpx9b_inst_0: DPX9B
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 9,
            BIT_WIDTH_1 => 9,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"B9DBADF63904B2E965B6D864174B4DCE4172B7DB2DF64905B6EB73B85A6416DB2DCADF4C",
            INIT_RAM_01 => X"B65B2CB73B0DA2A120975D2D36CB2C82CF6EB4D8EE769B85A6C961905CAEB74B2DD2C765",
            INIT_RAM_02 => X"39194C46936080E861101CCEA62349B8D266965CEEB74B2DB64173BADB2D965BA482E775",
            INIT_RAM_03 => X"3A9CCE069101CCEA73391D4C620329A4E873329B0DE6D100B0E865369844074349CC406F",
            INIT_RAM_04 => X"100804020399A4E86137194DC653B080E6693A9C4406D3A9B0EA62349D0E6652B0805C6D",
            INIT_RAM_05 => X"B85CEEB53904BAE969B65964173B7DCACB20B1D96DD20B1D96DD6FA24825D74B4DB2CB76",
            INIT_RAM_06 => X"B25A6C76EB4DD24173BADCED37290592D320B65CED36E9058ECB6E90596E773B4D92DD65",
            INIT_RAM_07 => X"39880E461371A4EC6C3A9C0406D309A4E845904824120904BAE56FB85B6CB74905D2DD75",
            INIT_RAM_08 => X"329C0E675298805C733A988D2633A984CC203A9944073349B0CA66101D0CA6D30880E869",
            INIT_RAM_09 => X"100B0E675361B0CA7410190DE6D399A4EA65101D0C2703A1D4D86F3B080CA73399A4C86E",
            INIT_RAM_0A => X"904BAE975905CEC374B9D96CF6590596EB67BAD864174B75D6C969B1DBAD3749058ECB6E",
            INIT_RAM_0B => X"B0DB2D975905D2EB2096586D96CBADBA4172B7DD2C775B0C82EB6590596EB71B9DA6EB51",
            INIT_RAM_0C => X"349CCD26E101CCEA6D349E0C26D101B4C24E904825D61B759EC36D905CACB70B95BEC76D",
            INIT_RAM_0D => X"381B4CA73101B4CA7310194E4653A9CCDE70101B8C273369D4C663308805863371D4DC20",
            INIT_RAM_0E => X"10080402010080E669361D4C66134880CA75389CCD275288805C733A9C0DA653A080E465",
            INIT_RAM_0F => X"BAC82E961B95964172B7DD2C775B0C82C969904B2DF74B9DD6D520B0DB2EB63B4DA2CB76",
            INIT_RAM_10 => X"BA586EB71B2DCEDD6FB1C82E775B6D86ED69AB4825D63B0C82E565B85CADF63B6D86D96C",
            INIT_RAM_11 => X"3A938402E399A4E669361A4C66133080C869905D6C772B0C82E769B65B2C376B75BEC720",
            INIT_RAM_12 => X"36080C274391BCE020369D4D875311A4E87332958402E349CCD26C3498CC26610184D86C",
            INIT_RAM_13 => X"399A4E669361A4C66133080E865369844074349CC402C309CCE66136880E865329C8DE61",
            INIT_RAM_14 => X"BAD8AD36EB4D9A4173B0DBACB63B2D869B20975D2C320B2DCAC36EB95BE4161B9DCEC36D",
            INIT_RAM_15 => X"A1C825D6DBADD2DD65B6DCACB6690586E574B2DCAC368B8482C96990586E773B0DB64173",
            INIT_RAM_16 => X"1018CC22031994DC6F220805C6D329C8DE6C90482C372B9596ED69BB482E961905CEC372",
            INIT_RAM_17 => X"10080402010080402010080402010080402010080402017194E86E30880E669381C8EA74",
            INIT_RAM_18 => X"100804020100804020100804020100804020100804020100804020100804020100804020",
            INIT_RAM_19 => X"904824120904824120904824120904824120904824120904824120904824120904824120",
            INIT_RAM_1A => X"904824120904824120904824120904824120904824120904824120904824120904824120",
            INIT_RAM_1B => X"3A9B84073349B0EA63309A44069311C8DE4D904824120904824120904824120904824120",
            INIT_RAM_1C => X"101B4C2693A114402E369D4E86334990406D3A9B0EA62349D0E6653B080C66110184D86C",
            INIT_RAM_1D => X"101CCCA63349C8E86C3A880DC69101CCD273349B0D26330998402C399BCE465101B4CA73",
            INIT_RAM_1E => X"B9D964165BADC6E769BAD46412EB65CED36E905D2CB67B2C82E769B65B2DF6D904B2E975",
            INIT_RAM_1F => X"B4D8EC36C904B2C320B9DA6D965B3482E961905D2CB65B95BEC36C904B2C36EB95D64174",
            INIT_RAM_20 => X"3A9944063329B8DE44100B8E46F3A1C8DE74904824120B6DD6C972B2DD2DD6990586D36E",
            INIT_RAM_21 => X"36984D86C3A880E675311A4C67530998402C399A4D86533080E861391944064379B4E669",
            INIT_RAM_22 => X"171D0CA6D30880E86939880DA75361D4C4693A1CCCA76101BCD26437880E465381C8DE63",
            INIT_RAM_23 => X"B4DC2E575BA482CB61BA5A6ED20B1D96DD6FA24825D78B2C82F165905CED375B8C82DD49",
            INIT_RAM_24 => X"BA5964161B4DBAD363B0DB24174B2DA6C972B2DC2DB6990596EB71B2DBA4163B2DBA4173",
            INIT_RAM_25 => X"329C8DE6C101D4CA2039984DC6531994C24D904824120904825D6DB0DA6C920B6596ED20",
            INIT_RAM_26 => X"321A44073349CCD26C3498CC266101D0C27538994E66E3798C406D309D4E22031984406D",
            INIT_RAM_27 => X"101D0C220309B0D87537080DC69101C8CA67329D0DC49100B8DE74399D4D42032194E620",
            INIT_RAM_28 => X"97586D96CBADBA4164B4C82DD69905CEEB74B1DD6D920BA596EB71B4DB2C320B2DD2DD61",
            INIT_RAM_29 => X"904824120904824120904824120904824120904824120904824120904824120904824120",
            INIT_RAM_2A => X"904824120904824120904824120904824120904824120904824120904824120904824120",
            INIT_RAM_2B => X"904824120904824120904824120904824120904824120904824120904824120904824120",
            INIT_RAM_2C => X"904824120904824120904824120904824120904824120904824120904824120904824120",
            INIT_RAM_2D => X"B9DBADF63904B2E965B6D864174B4DCE4172B7DB2DF64905B6EB73B85A6416DB2DCADF4C",
            INIT_RAM_2E => X"B9C82CB63B9DD68D20975D2D36CB2C82CF6EB4D8EE769B85A6C961905CAEB74B2DD2C765",
            INIT_RAM_2F => X"B75A6C975BA5A6C769B65B2DF73905BADF6E90586E972B7DC2412CB6DD6E770B4C82DB65",
            INIT_RAM_30 => X"B4D92DD65B85CEEB53904BADB69B7596416EB7DBA4173BADCEE575B1C825974B2D9ECB20",
            INIT_RAM_31 => X"90482E565B3D96E96EA4C825D6FB4D92DF20BA5A6E169B1DCEEB73905B2CB7690596E773",
            INIT_RAM_32 => X"B2DB2CB63B9C82E96EBAD92D363B75A6E920965A6EB6490586D975B1DA6D165BB482C969",
            INIT_RAM_33 => X"B65D6412CBA5A6D965BB482D973B4DBA4163B2DBADF44904BADB65B9C82CB75B8DCED372",
            INIT_RAM_34 => X"B6DD6C96EB2D8AD362904B2E775BA58EEB6C90482CB75B3DD6C320B0C82E765B1DA6E574",
            INIT_RAM_35 => X"905CEEB73B95D6C720B1DBAEB4E904BAE56FB65BEC920B2DD6E373B4DCACB6CB2D8EE720",
            INIT_RAM_36 => X"904824120B0DB2D975B7482CB75B3DBADF63905D2CB67B2C825969B1DCADF20B65CED36E",
            INIT_RAM_37 => X"B6DD6E96EB2DB6D364B75BEC720B6D86EB71B4DB28320975864172BADD2D363B4D9ACD65",
            INIT_RAM_38 => X"B95BEE16DB2DD24161904B2E96EBAD92D363B75A6E920B6D96E720B1D86416FB4D92DF20",
            INIT_RAM_39 => X"B9C82E973B2C82C765B7482DD61B2DBACB41904BAE961B4D9EEB65B3482E969B6596ED20",
            INIT_RAM_3A => X"905BADF6E90592CB53904BAE775B4DCAC376905CACB70B6D96E720BA5A6D965BB482C965",
            INIT_RAM_3B => X"904B2E975905D2E765905B6EB6CBAD8AD374B9D96ED20965CEEB62B4DBAD366905A6EB64",
            INIT_RAM_3C => X"904824120904824120904824120904824120904825D6DBADCEE169905B6C375B8DA6D961",
            INIT_RAM_3D => X"904824120904824120904824120904824120904824120904824120904824120904824120",
            INIT_RAM_3E => X"000000000000000000000000000000000000904824120904824120904824120904824120"
        )
        port map (
            DOA => dpx9b_inst_0_DOA_o,
            DOB => dpx9b_inst_0_DOB_o,
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpx9b_inst_0_BLKSELA_i,
            BLKSELB => dpx9b_inst_0_BLKSELB_i,
            ADA => dpx9b_inst_0_ADA_i,
            DIA => dpx9b_inst_0_DIA_i,
            ADB => dpx9b_inst_0_ADB_i,
            DIB => dpx9b_inst_0_DIB_i
        );

    dpx9b_inst_1: DPX9B
        generic map (
            READ_MODE0 => '0',
            READ_MODE1 => '0',
            WRITE_MODE0 => "00",
            WRITE_MODE1 => "00",
            BIT_WIDTH_0 => 9,
            BIT_WIDTH_1 => 9,
            RESET_MODE => "SYNC",
            BLK_SEL_0 => "000",
            BLK_SEL_1 => "000",
            INIT_RAM_00 => X"0381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E07",
            INIT_RAM_01 => X"0381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E07",
            INIT_RAM_02 => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0381C0E070381C0E070381C0E070381C0E07",
            INIT_RAM_03 => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F",
            INIT_RAM_04 => X"0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F",
            INIT_RAM_05 => X"0B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C16",
            INIT_RAM_06 => X"0B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C160B0582C16",
            INIT_RAM_07 => X"0F0783C1E0F0783C1E0F0783C1E0F0783C1E0B0582C160B0582C160B0582C160B0582C16",
            INIT_RAM_08 => X"0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
            INIT_RAM_09 => X"0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E",
            INIT_RAM_0A => X"128944A25128944A25128944A25128944A25128944A25128944A25128944A25128944A25",
            INIT_RAM_0B => X"128944A25128944A25128944A25128944A25128944A25128944A25128944A25128944A25",
            INIT_RAM_0C => X"168B45A2D168B45A2D168B45A2D168B45A2D128944A25128944A25128944A25128944A25",
            INIT_RAM_0D => X"168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D",
            INIT_RAM_0E => X"168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D",
            INIT_RAM_0F => X"1A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06834",
            INIT_RAM_10 => X"1A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D068341A0D06834",
            INIT_RAM_11 => X"1E0F0783C1E0F0783C1E0F0783C1E0F0783C1A0D068341A0D068341A0D068341A0D06834",
            INIT_RAM_12 => X"1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
            INIT_RAM_13 => X"1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C",
            INIT_RAM_14 => X"2190C86432190C86432190C86432190C86432190C86432190C86432190C86432190C8643",
            INIT_RAM_15 => X"2190C86432190C86432190C86432190C86432190C86432190C86432190C86432190C8643",
            INIT_RAM_16 => X"2592C964B2592C964B2592C964B2592C964B2190C86432190C86432190C86432190C8643",
            INIT_RAM_17 => X"2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B",
            INIT_RAM_18 => X"2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B2592C964B",
            INIT_RAM_19 => X"29148A45229148A45229148A45229148A45229148A45229148A45229148A45229148A452",
            INIT_RAM_1A => X"29148A45229148A45229148A45229148A45229148A45229148A45229148A45229148A452",
            INIT_RAM_1B => X"2D168B45A2D168B45A2D168B45A2D168B45A29148A45229148A45229148A45229148A452",
            INIT_RAM_1C => X"2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A",
            INIT_RAM_1D => X"2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A2D168B45A",
            INIT_RAM_1E => X"30984C26130984C26130984C26130984C26130984C26130984C26130984C26130984C261",
            INIT_RAM_1F => X"30984C26130984C26130984C26130984C26130984C26130984C26130984C26130984C261",
            INIT_RAM_20 => X"349A4D269349A4D269349A4D269349A4D26930984C26130984C26130984C26130984C261",
            INIT_RAM_21 => X"349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269",
            INIT_RAM_22 => X"349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269349A4D269",
            INIT_RAM_23 => X"381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070",
            INIT_RAM_24 => X"381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070381C0E070",
            INIT_RAM_25 => X"3C1E0F0783C1E0F0783C1E0F0783C1E0F078381C0E070381C0E070381C0E070381C0E070",
            INIT_RAM_26 => X"3C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F078",
            INIT_RAM_27 => X"3C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F078",
            INIT_RAM_28 => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_29 => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_2A => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_2B => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_2C => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_2D => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_2E => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_2F => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_30 => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_31 => X"43A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E8743A1D0E87",
            INIT_RAM_32 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_33 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_34 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_35 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_36 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_37 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_38 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_39 => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_3A => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_3B => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_3C => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_3D => X"83C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F0783C1E0F07",
            INIT_RAM_3E => X"00000000000000000000000000000000000083C1E0F0783C1E0F0783C1E0F0783C1E0F07"
        )
        port map (
            DOA => dpx9b_inst_1_DOA_o,
            DOB => dpx9b_inst_1_DOB_o,
            CLKA => clka,
            OCEA => ocea,
            CEA => cea,
            RESETA => reseta,
            WREA => wrea,
            CLKB => clkb,
            OCEB => oceb,
            CEB => ceb,
            RESETB => resetb,
            WREB => wreb,
            BLKSELA => dpx9b_inst_1_BLKSELA_i,
            BLKSELB => dpx9b_inst_1_BLKSELB_i,
            ADA => dpx9b_inst_1_ADA_i,
            DIA => dpx9b_inst_1_DIA_i,
            ADB => dpx9b_inst_1_ADB_i,
            DIB => dpx9b_inst_1_DIB_i
        );

end Behavioral; --vga_sample_buf
