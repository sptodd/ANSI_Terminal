--
--Written by GowinSynthesis
--Tool Version "V1.9.10.03 (64-bit)"
--Fri Nov  8 11:09:02 2024

--Source file index table:
--file0 "\C:/Gowin/Gowin_V1.9.10.03_x64/IDE/ipcore/DVI_TX/data/dvi_tx_top.v"
--file1 "\C:/Gowin/Gowin_V1.9.10.03_x64/IDE/ipcore/DVI_TX/data/rgb2dvi.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
ReOVIvgxOP1KC3oxLReiFakuTn8OYyhjuLfIJtzEhfUEMHNUSDGU5Lj+5ra48TP01x6HnoCg4E4a
K6iJxtZWSidgxznXrtquEecmrIR+x9yx6bY7HD1xM9M3kZ4Oiwo3WMw8IFXQ9ZpvKTiLGm5j3bTQ
WjI44iVRElWaAVxGDrmCFoWwndDKB54nDyPYRLdg5Nlzg7WyrJg0DC2KM8nK5b/c+kGVLZfb6Pi/
JQjrMOZgw25bXaWeNF2NTeND4O3If7+9os0wPbRfLDbS9m0u7oogCnkHsTJDOnKeQvINLA1it5Ff
F1gPaM5giNkboBUFaxF2z8FUUQPskSthxyZw3g==

`protect encoding=(enctype="base64", line_length=76, bytes=67200)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
mpyxUkSj1IMcEeGXdoJWG30KPr68sTLq/xLzzT+kZQJwdqCnEXFnoajasPS9vBozKj/5uOqJfkgy
fQKEMjOccQrk0cOpxoLYMHYfkgc6kiHQUd4WaA5B4n92F6xv8R0sxZi/cjP/pHK20YBPaoUXEJIg
1qnNfaO8AREgpn8SEeBmM5dJuClHp5Ja+Ldk054vh5KyUNnDCCu1tfvvRtLi7ZxKRyTQBYwM2Y8s
mzcPKHVHwTifx2qP7AFeJD6kQAlfOlFpKkbpuce/Z7ELP1Di3iqlW54RWlO2MRm+Cgd6EdDLFKyn
fGVWJwRO5E5BNh+uuRTWvV/8kZHxxu+gPlSJkhfHAXzD7fuMr6oLjKHPGbwerU//vpwyoWIUKN9r
qUjXOaYuIA2batsNvsd8A7G2nwQ592eLQO5UHfAP8NnPIUxuRBg5oBOVKhtQ83VrKn2+0S8Vfw/P
5K/iNlouOxhbTmVTf2uvVdQU3EmE6S73aoPuta7AMiT5d/V2bVxPXSZ4u9/MuLN/TILMmWebsHNG
V5PE8/7A4gGcLwIbC3wTMLukxa66mmrUGBebOTMZ2ub2Px8fNXSwQH0cM4BVAUzlgxfiP/x87NF+
ewNfgMqoTp9pr3cIT6lzS6eK+MIFEIfHXn2Fuigg50yRrb1/Z122OuZGq9/GzAuVg7S7se2KREj2
uTYCq+LnCW84KkUBVoIOby+9Kkc6dcdMuwWEguP5tY1MHo+EiR3IiMOQpPo+x/e1HA7Dwh51OmB9
MuatZUlboynhBH7BvXB5zMoIHgtVGz2sHeuQLw8aazFHVAAesyslFfgY4ZoKd4evDgn3Wm3fGauY
7zhaCM8Jb/qyfHMTS58EcqHMu+ra8JCR42zov/gS0tVfqzFK/tiOxKUlgAB5Vq1n+2WleTyl3Vm6
+NvJVCSeYX8fzl2kA0cgF+coml1R5JzEtbugJ+GoECUypgafedOh2SDX+THEvftM31jBWWT+wpXL
wV0qhv8RzmEf/oyfB5sFJ1ZtRSZfXpDw70vGOZsDCao+UoTW6dUO0KMY3QgUPCmziFHwbhtOU7KN
V8FwKQSYlt1/PAPC6sjxnFr63kZ78yGcM0YbbGWU9lWyNwreXXKz50YSFM4hmxUZldqCSfyqO+D2
Bvd5kEpNo0hSxK/nUUJjC8PUfzmGFadhxxjUjAbXQs39iT8EJSQLIMgpzOmfLm4l3z02x3eM8cX3
il9q/pUe8LmSttpxxHPtJpgwzTGn19yU4UWS6n7A9rC3fy6QHEA1m9eSbHi/y74Y1jChYRSjOBjU
UJjZ6m5uHpQfvzoTuYP/7F1PzB+DoiKx+blYrGZf2nvEYy+y0wTir1R/hewpEzbAyXg5ASqacmn7
dzzq7+1xzVMAK9XB2AKH7twatiwwLbL1PSsral7uZ22p97S+VJnA+CryORH8u4oVKkgvz2pkI1sG
mRd+xesZtLR7JSkIqZ1q/FSAfCFoEmcpKfDr422Xa1SOfuqI/+3qbfM0H8QKmT+AHJv3s461T9eQ
t0KvBqDFZBDf4GoVzHINMc+2cTVjCYgDOa5ZFGmcihmhB3j9sNZpGhnNXCVvX49IkbCartUmru2F
bqPhZufDxfO5LSDtdAOl3Qn1n5A1MlcdSqJE0TlzyjQ3XHSD8mP1z7HKBsKYIHfGpreY7caiCRI4
cDB6zC3eqQ0mLY7YURpQBvIaK4xRHRz63tojCkqNFTCNrIz8qa2ziea/sBhCD1dPyHU5p00LFkEb
OyPLrdGYOvQCRxzO70Q5TZdR/fAFNOLPB6+8sqLUin5A6p0bez+ry0i/XzjtAXrBp/kI+TuzdgG4
d8M1bJfygQ8DjuSmTl+cTpK0fCchiHtGKbJuxe5UrEPMvHou9KzbGPw8qx0kRpV/BstB7I5M4OuD
pR/fBgjxDlecgQT0DQeeG197mZIZCKjoV3cqV0C/fnXOuG1pghGAJTCUl0VdQEVX/A8V/FmfLGj3
zD99CV1ZBjmhzthy6HDxeFVwp2Iye0hTaqdXpzSskHFfs1CRB9ea7UcL7uEVeD7ozGbnvOKgqOst
pJdntd1mdf2mBo17p9NsB8ANtWSqUzZA88Razpryy2YL/W5MJsRu1UyK58d13oSPC4EkCscA1XBQ
USRC0X4h/gRadrY3Lt2Gk0j6C6dpQov0JVdy8e3yTyjnvV9oFcpduqk+LIW0abowFz0vAN58Eq81
S6mGQO7gkTOGJKW+ZyUSpLUJSaHkpxS2SmMXVIX+BKXCXPcD5TN4wejygLDpqGRhNXMoLZyeTr8S
3XgmakYXZ6XMTfCoIgb6wNBJkafqOYGQaah5VJk9cyeOv6DnWgfGreMvQ5SnpcYYM5JOy65fDOmf
Id/JM05oMgEQyeErLGxqXLqMEddtDQGxjcR+HEu8ltUyvjZg06n+lzzvav5sa4OSVsP6QM7qUq5O
rXtMk0JU+dHwLrPNVT2CIYY4/3kDkUU9/JnRycokECqh2ZRTKP/lbSdT4h+FuzHyHVhqkdMyhr4v
LdhZ6kq6EfZR0wGrOy81f73eLXf9h7EIjWCKzkvoocKS1BYVt/wtpfegcCYOvaaZtzKrVCRn3fcS
MjxsClUHwSTkhYyeYme2fY5twvkQh669jcV86RbRrJdfqbewI22KzRl/g9XhlfNRIp8e/PjcGuVQ
7HWS+8Pcu1+TIKXUIzVZ+U3Ed6NP9ZD0Ziu1sH5w04DUvmo00YJT9VgKeSILpJZi4t2tT2Vzj9o7
+kSHWVWKp5U7DKWOvBhSD7hdyxX9oOxDUOpjtve2N4WpaK5zT5B8Z/VVfDubnl4GMBZxD8jJDpQj
8J0sG9qqJoGOrteWahBlb7X3h4062a/rAmbA7hW7y9V115DevvjA3xeyV1LoBeqGqFcN7UI0vycl
cjijKS53y9qQB4Eeu3ip5pOa5L6T/LEXoZiic/Dm6/KeLIcW4y2+880xrvBEEVvxR/cUKQdaoPCu
omp5cXFgg4z/lY72hK0iX2MPKpw3UzgGJik/MCO/8+RVwMq9qNwOhwipwfy/FJAAoV2UC5GU2FSs
gM00LQwa1uz6tvQgcaVzLhoIFARzCbFy7hIB1r8ZvSZ1vYm7jUmKFwFOmsUcDRcsSKiVJOeG3ViL
TfgLcnTYriQ29fK67KcgiOtZcvvBbhG73nnwe0Wbmh5GLvCSqvMyXumfzZH43cFFRekpvv+35lI8
KEq9kJou92oq45SUqoJfTmZ5l5PN06hfTCOll9ywCd4NPhPAW9QbFz02da3w/QrM14kJXWE6Zbkn
uVkjYSTiRX1SK4OaoYGOsKLBXsZ2hAp549Xr5GeELov4Y7XiyBlxgAIk6MFApEhNhIS3y2P6qoCS
7q9M4NOvhJaDp2vLybxc8O0fFyiyw9rPsxRmTqKpeUu+bbx3mvLpyKRDLiE6GGN32fTWF5rsA4z4
6MnU2SERguaDck/3AFZa+BP5Nrl5VkYnCB3qyPhA694LGqvWv6L/rcz+oBK2v+yz5Y0TcbZGk6xo
P0Cl1SMcAS2p5/gzVGjZNf7yiKuqFhbxHBZ9yuwHs733tf2lr7kiLOP7LJgbcwBYFV+1GNXNVEOg
IuZ39ChnUpzr///H14Jczf/2YQHWVeqE2OXvIldyElr00ViaIwse4VIsNg/niTUy4dRH0JRIfiWA
cv4m0UxstUuHHgnxdDKzk2dr5+M8LgcnrKfPqQfR4m/7wmNrk8GfqrLs5Yl/6xb/u6RCuswZe4xN
pA/Bslk0saDdvurm+2ahj6fge5dYmrYla/Eu7Xpw9XrgsS1rH8ySp5rDyEST2k3doSY1mj47P2Le
hXH8TpmAUVLQJvFuhuKWL1vxpX7hwnusl+cbphoozCZzBlB88u4NSOVv3yNbjNxmW993koZ9fhMp
GSi7XdHTQfeGbsTV7olGoDGn0p8BTHhtbNm7so0W1ak6rf6pooS7RbihicfeXRNzSuhl1quP1uO7
FeqTnAVY708vreehyCFB+bTkH4iHt9DfPRv4/snvkU5/WJH7fsYkQhbieeZ6OHGl5627Uh8PglRC
htrjkczUaLmKS6JMjmS3TImcXT1+uzbKSbbBM4Xye22NLI3XOw157OJNJ7QZdT/+tbboq76WnRIb
bkleri/akAGLBjhSZTUYBLUH9FU9RUlmeNK48KmH0bTdPwQHRhMncP2ll0Fa5pA0IvXSUVt0Pcw8
Yw1voEL2lRFsPm+n/glxivyMzpZC0RVsvqDu6PpjdV5UU3U1mGU/9P+v3sxerfvVcV0B5E3mBMXc
KokaH4x4sTBzoABE3L8f/sX6Qgd46h5Ker5Jyu1rEVqOFpheCcK6d/+bsKuN4DWCt0guZ71p5xLC
il/xGbQjaaxg6AA0/hX70mUsqp7bpL/egWrsShBuTKGnaOzTjCGCkk6QosYhdkajDsnV49CdU3m9
YzCvlGs4zu86CgRBESIZ1WipvQwlsFRIsLQIX7gcvQ74qrcGAYiUzhpDntBmnZluvlRziGZZaawg
EqTBD0hTnejGIoRosChbkiat37E7/8NjQ+N73E2pkai9nzNrNk2NUYbismf91CXhhHnCll1ofrem
Gnsr/7tsvuqvj5k2TxmGE+whBhlAQqBwD5fAet1N0gDWqWyb9S2KP+pR+D1NhU13Z27Z6hIkB6Nz
ieUNPiSt6qYXc/Z7cvXZKXDU6quRscNUFHzG7sQwatShJO7BIVmrGZI7ivmsCYHssb55+LA7/e7n
A9QnlDybS+N5CVDtBOa9PicDATnv+m+QKjfHKsGxYbMVBgnEJ1ta8VKSBYCYZLSzYxPK0oJ9V5VU
BdRvp0AvFNuatB2rjZGsIaBc56mOCiF5vP6qiFdMM0lVu6dSg5EYV8S+jXWYkK4Lbz2+PZPrdzHE
PqdxrNnrGny53SkW12X5c8pM6XYNxmto7s7CFRJR7rpI2rZBCuYs77SKrYqfcuFJ4W89AMkSAwm8
0wroa11haSYAB2d8rxdYrkB/6hS3gr9K3WtsRxBM+me+mA2S/kmso6MfmYLgu4tv1P3g7er+i9gz
x61Yvt2nb8U0rbynyXcWHupZCy13Tzu2jUKzbwobI9SzM1pBl8jt8Ae7X5C0pDmau7ebNMa7fy+D
U4Zl3WzZz6zBOkyW3o/EXQjA6T1jIwvlj2BCDwJxV0GiaDVZleOJ6oghbxKmrhgW8m6xEj25zbxf
GpQnoIZfD1r51u5I6Lv1sGpvpfQSCRGyRq3xwwscZfXCvBePSi+N0tEH+dZOxj+wSp4OK7Z8PkQL
H8LqOlgzf1hMljj1q6b17ddljY1eV+052brYeQGluhko/iWwn1TRtzx1FE102rcbjh8v37hn6kpV
tqR+MRkiDKo+WURqBfAiumHTIqxqcpWUkNynYIfCITtsQ/iqn3EhxnpOOAl2hFBulb8TU9/dWHwc
6xgYJtuRh0zZ71EL6TxXudC1K0kXLeRyrcQK6ARBcKqFoLR/nkZBXkJPKtHR7dXfFToOwWhjYIq4
drb+3rk1bhlGdW4YQRMRQJxHp3JuL/6vWDs3T49cLg4Hq//OWIAZayUVQQQL+ZlWZHJYWbHnSeXq
gnw66dzIQ4JB7teBo/u2ln4tnyum/OPt6+LB/fTb8kmaNt30fnlSD2f/WkL2E/3yCgaOrLPpYN1w
ls03dNCndqGsfxjJa/suBFtKHlEEu8aZ4q31etQuv98INr8GOdK6ny3p33M5+IfLcGhG2gAfj+Az
HIH0IVJ4SPpd0npgEsnj8rlfJmUNIaykLNmlZAnaFZvdybrROBywRArYdSmmgnNFYy8WfY/Nde2d
o2JLEDRFlRlkY7JG9IoqtJZy8gCmL5sY7RyulS6y4Zb/G8sHEvCzu2IMCBb4iAS5f6YXrj3boZVT
pOSRFWVoz9oz7VkyRIbjPIAet3ko3g1oAHgfkenIql1AYAqSrfaJB1g1ECIyAn7o8L7g6Yn2XjIM
/FM3zFzILLg32fmsfjSGt2JH/UwkDQ4GzPd/IS2juMPCtJf3aw8snWe9ks4nd7wTHnphtIbqDb5Y
hN2c1hE/cFln4qHGcsebDnV474tdQ9seHwCk64tu8uDCHRb91mPbXLoa2h5vpt07Vb1qg5s3APaq
hguyUdXINPafHdMTDlRENRdZS8SOdk4YmPq5h0aF0fwbDrY5IaLPk6eYYY3UcHGp5/605vattZER
B2GhTle24uSKrcSXacuB+uJLNXov8Lx0K1uJDprSHJypJW9qOT6TdMWr94oNe3EW4taLT4joG9Ll
5DEpQ7SoFRPF13dWGmD2YgBpl3PZnRRjVsRoE1izHli3irA07Jv2/RSY9TL/0KrFC4WMBRsgvTN6
j1aXh1mwKMmplTLxP6lRnIwiWz6N8b/J5yUiaiCv5ouT1SP2l+b0kIFvFdVkyfKqOB3zTCIBBYod
+9rQvjxvNC4Gbg8UHEr4iPyMLk3P1Pgic3+tWzWxI+FAIirlM3Ngz3xLl3GANggCHkw5F7GNRQ2X
QSwMdqHQpft761YW0ccTM1Uxg8wdb9W9RTGOYVP4Foezo/UgXW88pS6l5kgBglWlvUluqDzHGZNX
GMu1LsT0Jv9JU43xB1efPwGoSHAw827LLMHOwys14VYzvSxENpCTHAHoAet1OigrXHx4EuYln3YO
K2ZhMRNakwElqIp0j17dESZ8WULbjHel2DwJsg8LS14HfVlS0iWtL8rXyvChrWu60210gf/PTb3J
JbJ7MCYqdujuF9jh6hpQjZYr7OWQKsXHYdqBiUMGJUFpcbPJyzruWwiXkfOIfv++EuYNX8qsG927
LBZO14V77ZdKBbypHmbgaJnBH1TFFl/QCLsYquz1S2TlgMO+E7HlpxzbrjPxeLQfwRMFFZw9Phhz
3Ff8HTeu3787YZwLwyL8HDPCmNV+pwotzFDJ2wnCgt4OTizYrYfNGF/gEartkwAuvqNBXxY8wKaT
fw+va9DJH/AXqS+syN2MD8QqeHBmBqqQ+HZmf5YNiuG7Kgt/COjnxLLVQkkBErjGy30WK9SuF13x
na1ok8xTea8NqujYm2BnzbQHI7C1gTGT748TptqAOf2IPwicgPlY6DbC0y+opniEK8dof5V6IyBt
1MxHGv2ysAYe77t1CT2Zt9fpx1lyRr6NNmzTeEpnSYg3yqBukQ1EPtAPsQ0lXnE1JGB3DYJVfcN9
Qf/U29ZjmMS9km24AeeYHoLrDClwY5eOoxQ3Zz1pNk4lz5XQu/GBEO3KGIihzcF3rfWJ911FzjkJ
BZ/IsXbt/sYbGMLrGz9F6MhzqS8njU0e56APsGcQi9/p0xCxJhwg5vRyaqFG3NIioZRPvTfGAXev
XYV6Mt/VVcU8iH742W9YWkYybJDWJwaD7grbw1wx4udPMARYbGKrBi4Qm3S7Hww0ApH0xDVign+z
EG/Cp2nX18l4WMUeUnees+72XIpfl3u3MNmRrQe27nu+5Evwue6ZCO6RDhaUICmDyNmI01oxfpDI
wfZmz3h2hizZMa+PiagYJ2QlHIHCF2a2ClxvVS1N/j7T6S0KQ0lZ+fk00Yk+YRJpL7EXTnMl8H2q
1K5R35GtWO/8wcPSJ4275Oc+CcrYGMTssISWYfOkE1pbza6+x21EJFkUAmdNZcfzofp3pjlieQos
UbiNfTZ+FgmgCVxv1ctwmvgDMElNaYQLR0+hEXu7MKnfYHYgabiMp/pF5YfXF6j1EPeOzeZxduX6
cKtWW7cWSY/MkK9zxdEK31t/4TQKuICQwXOKN5d13mgGe+sWppE2rsM5NkdI7Iry3AepiI+btBpR
KHioHOvKtDJW9rS79A9eP1R+WEtsCujgrg53pYRu9GfzxQTgkz4kKRkk8ePYXu3ZmqHYB6h/Zpbl
ZlIUHt2f94QLTaWEm2qzMfRPOOEhoIJ46DxS8d6e+hAzHPZDNef2MGhWvpOuRupFDR1nVsNq86Yp
xcNBUyU+VH1ZVH/sEOPA1KFQBS/dDw0kuFmt26hvOq6ciUiG30dV7w6ECyjbI/P47cnoLS8NGqqj
loCAM31LBvU7Jojm9HBiGu/ObaOpUlLYUtySADw/8g4atKKQv5pRtCeJeXZMeGJhJtFqxNxHbLkp
oQbG28z93khZ4Ek6u9T8+vd74Fg0IZVHOZqwPMDHwnwmptFINrnWIvkuxnyMOwJi30+tjp0cXomW
4p08AtAZs8XaB6nP8b+u72JyA9WOSA2Two2Hx0+Ii7il8fbKOls9ux8L8+qy11QXlFUiWQEYygqJ
JvnvdO9Q39xoUftCOuC5ZQsuN6cmCHsoBbrMQnDCmIbyU7nG4xBZkQRK+j+Kvxqx+rODvT0tmEe5
eG/RDTALD+/PftwAhep3hTyZbeobrwwQ8Qq1OO3EPSxLJ3pwdFG1BB3eUiCoHLXN6sbahPuWJ5yk
rP51khTlfA7QlqzuApYlS28Ym//yXBOll7NRTOOwSerLFROAUIc8bjLc7ZS9abByLrwObmKoRTik
akIDauzA6X+757tCSkSzOcC3pmhcYmavw/SulqBQ6lI/ELzHzmNs291IqQdJJiEQsu3kTdOqF8qx
piwhNJzwRnT+2bflUKsqDSYpiDXPIDEHhMgKLayVs8zLXiKN5azwdAVJCfFnCt3Y+TYhQbXLHGBQ
qSTf763VtjkUMNBz8u1MOk4P0AR1ddIJjfjZt8Oxe1khfUZUQEp9b6nt88vzQaL60wFxPty1NdiO
E5B6jb8LZBJjJLhMmZrXmzwmiACKIasWCycQfEZS2CJgIc4Pvtgqiy/Afr7mg6xMy6MaEEEaCAhK
5jqqf8jA9bZu6WFz3DigyIbvf+GvGEHh5WGnlAclRAkOB6WNGk7KkdmmTkO0mQjRLn5XJ0ZWAxkU
I4mnwmk5xt/wORgmZH9mLKtprkTJu+lkkXL1ivbEGRbY0JEoKIWWUMaIBjgMNi22g0rcGHM7N1pY
xy29RTDsavNB/VpKXqzo9wjtfJct/ItVYDLznDYeJoFJ53lJAL3bAaCDRF769ky3VuUaQA+X5N/I
j4bvIK41na+WKap2YhJAcOCx8BKHwsJeetjFN9OJeyaAT7C3Jwwznbb52WUOnsrnU3vDiQX92jVM
K34gYK0XmvQeWK54P66tQLU8vFES52kOpMSWn54eyGmHAB1KJ+wycaJLbF88a3nqUthpWO9kXSc7
+2WRc27TNsBuTfkLH7kdJCGBgYD396biYTLvG8hMNUcfz9vGwfn3l0HFbbFUYVIwFZmmpUjFRhAp
cV3TukkY0FdUrp2H+LRpyIjFHJnTu05PFYmj3b4O+YOWvuruZEgrmkvv7k3lE/5m6WBV0N4X/c2v
E2ynxcU3aTtsx/DPH6BSnoCGK453lV6aQYXaf3DKUgJJjtm6Hyw1OnoAICcDxP2F42Wdwfm72mpM
AGXe6ctPMJiyUr+RtdnULlX9Itas5OQJLd3+1UaOnMJHbu+KFTsnxfgy2iGamyB/JBkFU3h9tg+y
y66B07h4jQbYdGk2T5xqp7/qinpCaAMWmA+dtTIugig9eIZdV8ew/FPfNrk+TyeOtB2TVTUNHC/q
NRA+YIOXwQHDf3GXQQpg5119sC1BbSBhIGqlfmTsbdN5vEv1kce5i8t6QaJ5syA8V8k/6NnvypL7
QvlCfhIsuCthDVQ55e8Rh4Z36Z/9QqvI9wLETL0PZ4f1vZ9OcP3wX37nFQ2Fq9ZTyuJpyoGjvfyX
1V8zRI5dE8foFE8WRfYzLsgKKq7poXycxm9NA4UEIMwujS1mYeEe9ANkmOTNHcDsFb5Jcu6CjSR9
msfiyYGyCbO0HMNqwgVJ45ps2n1k+wDPKBKtM0lHc9PFQluNbx7jDuc4Uc1zp9EhvDTFIgmUsUNX
HJI8i49SJ608PZYOlPVaZaL58IgywQccIWSyiy8cjsWjozoHk3CZx7xSn8tYgnY8KjSMcp9+sEdX
LJCA0TpM9Mzzi8SQpfd/KR5sexSWMz6olZHpsWbZ3LbbYxkx/XZcjlgzFbMMskX69Xdw5W0mwDGi
eGAwaB/1izOoeR7LAIa1qOcih5heVMi0SFWNJL5VhYzwxlnyZRcEwTGYPhSQekqa82mkxQrZ45eg
KzYBj+3hMUHRJk8C7yFA/Wh0NIjEOuIG+vGlfGfObOaNP8LtyxENNAYHwKHmPZpFjpW5LZWnUNGd
1XQpPzicAGqdRx3ut+jeJ9ifbYqmvnwNXl3a40GKKNCsqFQURDOQWvosYFN3bIHAFLNSC3f1SFFz
bwWSDJKvXyvTShwk08PPbJU3lEoEYsmU+48w8YJt5RxgsQl0OHmIGUbWKG2KrApQSmUv3FoiXUok
WJ96DqQRxbhzDrUO3frjMyFePCb4t6m+lRzbSBtorTzcriZD51HNI0FaaD1gS4D3DgMjxtT3NHkp
S11TOXvaKuBbB63i2BwQ5pbypaHxHYeXjP8D55z1aDpUbxkdDRIBP8abM64S/NaiyibBCmsq5WnM
5/MSINyjAQ6SWUZAqFj9FoknX8XBXlnvYD5dBAAPSOY0oAg754jNRJevFNrmZthxz2P0kOXvZg0W
vEPeED+ACuSVitsRFg3Lo1mk34TlC9QD2Du+OSZ20O4Wl2cxMiBl3Z6LE8nA0U/qrknAXQ1E7LUd
2uD3vXC8OOKqhDXb/18II/drRhG1iyr4EL8qG7hWO/P9e4f2SaaMWXZ7hRiwzngsI1pV55Z8xMGZ
0P75p31peTgEChsQp/7Ol+MRYnwAfWyla/ckiZT3g9V3UlDY2bSixjOdNDXOvCzftZ2inWMRcdab
92PGLa7hmeCKonAhsmwrnmFV8XlCaACDTmW8seD0MlgGWJ5uLUw9P8UAvU43N9UvXyQirmr8iULF
cX3XGLucEZrLeqE72xtI/QsMKuXY2tnbkf4bVnY/f+4dt1mVVZPe9qbkeseoeMM1zmI5cQxFtSP6
X92V6qlkuiOqfLkUtEiN4wCsnfDlfwPVCjqYafilHscPxOrfSZuFJDc5T4dva96BojqJGyuYd0zy
N1jkslcbLGlRHPJdOlLU1TUPo1AOD/L930uKXA9bXvhWqSgYsi6Md/DUpRyXJBrGVvmbCZlYc2wh
54ueMv+TVMsprwzxlKSQDrTw5X2Pa7LqFB7Mn81lI1EIEgeuYogG1Rv4BdqXwrq394v2TFnEOU0N
ZkpWSuVXF9WeLS4YM7Vx0Qh+1zpH5ZBlrnWyXq7WllCefh+VKfetZPNIaWlWC4D5jxfrJGCRwdcO
yemY+CJUdVckvI8/jBGp0b+bqqdwcXKzekqPfL/GfQUzhBKM4Jmm6ADRsDe81y8RE8XLLtEb24An
Cb9A5LxLHqNaH4ga6jF9FI+wwkN6dG2ACzvi9WmW7xaq/akBGvaNJ/6+oEJnnUZK8GkqgbEcUaLH
wNfTj9N1gg2wrzLDpAZgOFkiPx04v2dbiaOAqawpq0eO76Qo15XL2y2QW7HSjUCKK2jqHIpQ2t9x
ZwOm3UK1af5kU2K8vPdyGUon89rjRpEW3+rNurrFvczGkgWPk9o/9XNbIU9CkVFuF5VhJU4cTT5C
tC0uWwSMkWv7gqxlzbxztJHYX2ivOEzeh/MDO+gz8qOE2Ee49kkI4w2j/DbszYtm1/DXSJq8Zl2h
km/CHrBo2PCzNF/acHalt2qiRHXZAnBPy53q/iauXqI19UfiEfIWuFrjyyeQHgdN389qEzavFSA7
TFzX++lWPOJa/bmvIUfFhZwCSSP2juOIef4tIKLeOamSEzb7uYI3QSVcQvcQ82o2ahkamVz8YuOe
Z89vWcXrpK8DtzUrsempc5UmSlOyQlQeeFS+pzrhuRNZeH8ZkbAi9jXS53Nwr2x4B7GtO943cGlB
+AodtFvN1I1MRxp8vGe/jRuC5TSuTElJB1+6lfeV6WUwMiWxLYn7XfGxy499HU+Pfg6GDn1XeXBt
5OHdwV52u16weKOfLI3u4a7pVWHHYZTJwWD6+5AnPFJQr7cGMDxzP9ZQG4HRbu+7Xtge4AxHx/M9
CdbvVkBYIYyewxJk0xwAhTtoKG4SUTyDBpvU1BvBZhPs3KCBEEEgmR9m/Sp4ZidTnAOwLtuJRH3W
iwxv6f3GX77hXmOfdHJhAWSBtLa/H1NjFadNu06Yk5tR4vu4eiab4yv+VEAqmd0VGTTJD07yPZHK
q4OWcaVPoDCULZP47VsKQm2j8REBE8J0eANYd0dePkPnfJf5YZ2d/ztNlt0/7NtGP7wacIj+y0sk
AXCHTKQV2SPDI8PFKFk+rEN1PIs8eIvHAEU8TE+n0QGMSehtgChdjOU3D6ZifPeJCKb3txiwXJUC
HP9IphLrOdA18Q+iELC+wzgtFZhhnFUPDpZ1TxOgwY32fZkDI7N8BGvK+tRgJnutPOx29LhVxbwh
hS48t03/OZfFTMiYyYdgYcnMtsQiU0TJAFjSRremjWQez8ehQeaRdtyy3W1ssGXcPav8FiBsb2nC
JAAB6LwtcknzqXJVpEraqqBTI4XGQb0003iYqxH2/jLaDsgmlOy7sbJ2C9maVDAhPA7O+ujPnU0p
9dzHTRwzG39ZVmFgXnktpkkMHB5jz9F/6EroYlFKCLQqCV5xwEjbpWbBe39GoGLzoikgFZPfmCCE
xsRTmBbRFYDECvhg4TLgiFMo/V2R0KDzk3zaJJ5eLnxtl4D8JFlIHTtJ7Wwby7bqJciosdo6yjJR
lcGUq0SbCKLjHSB+eOcGY9EUjW8abLprlr6cNkTiGBTGqI9G7Uz+hUIcvqw3PXed5ya30F/4F5K2
en4B4mppZSMiaSl40XSkMaJIw/SFMqD6t+vxUFaFyfReShYRkg/K4ZTs1M1eKC2o3Kwur84KnX2M
IBFcO+rfOJmZNawS+bNV3EpCZudIjXdwqT4oofOmZLe1bXiOuf/+MuP3+vrP0oT/F5luX99hyqMS
g4zGy0C2whEQLeKr3bRCoVdA+Bwn0ANVOnI4d8oGY+AQI6P+Dj9KRcbqPjWGnxQ8sT7sAJfmBkGC
Z7OxeOBiBjiyIGGzeHeaz5XDfPdFHpxjz11zzq+CkZXtYDWEQykjWscVQzW8bWainR50+2WXqVwA
9SQ9IqgmLA9ylNjpC1bZHbacXEJbEtoFxk9Rf051/cOrXcqpWgVaAAuhEVS4rbXX+LAksMwdcPmH
9u7tLMuxQXv0IQRILssCHqutf4T+5ZtQEKo/0AuXeeLXkFeRtAkXTzGbxbVD5YbIjpYs+UzlNzHI
Brz5eZy1G1zZGUP4OcAuUDHw4yqq1k8ygg/aDEPonfkAy41JFqIRYwLU2B9/9aDEvBeq3A1aI8Dv
0OkKSNes9gPnbiE1ukG5AiQkPb/RlRw2LAblj5lEO7ci7DqArQ3MPFOccDDJxl89mXmF8jXkw0+f
kBzqieE8M0sIyOhB4H0P5fTmVQv2CE/T1qaDnyng0lLhbx6B6T8Y2dR4ByBHoGBA7ySBQY5CDFYp
Qv0JnbxKk8Bd4Aofkv5TX95ywdFYpdw/MYUY50qNqxbVi4Nu5DIyLIfnfECq24OdT3FFtmbmnnvV
PqIgNDTbixfymr7RXwe/a5qRmL0pzITwl+JoGDMKS8EL6ZkfBrpyDJYZ8m+HaJDtm/pDANSGXkTR
NUxQrCQjIEELqMNfrLgcfzQlSrfMdvDOSnUI/MI7o7ItCAd0zdACKpeF0mNh36rzGO9GuXc8ucAm
bxQbjyB+ofbQmLr6ARclwHMJAphOQiTVqmHC/R4K3zG+EXZn0GcNGTIbEdkDc3X/CMlWijpCUF5/
JEIDpx8y2RWK+LfcDTFN9a5GVFvHSh9wu5xBhYJgCIkmjC193KycUI21n98cb1DbnDrihr4e046z
NezEcwTtF9blekJ5HPRJSoZXkc3CZox47UWbt4CwIexQJy5ull49qG6/6MjMmIQfSQMXRIgdNRvp
0udzkQb6dUX/Lkyy71fjX96T4FZrf8N/EACem79SzM8qnfVqJmf9Neq3A9UteC4ojqToRTiNWY9P
adaZDE5jSDpCJtPST/yxA8tL/eQYvu8u2UJ3axaizxTDYynOmnzr4B0wLlm5D4R7Qjdg67OAI7Ty
lu4q15qbEUZ9PVwKX+coszxqc7XwBCUPT/YpIA1UBTVHwzmt6vYCMXZs1v0TixWQAAKWvzEu+SXo
9j8wiIZlS3QB6IkXuMw4HqZn8QgiNQknXU+GCe4tYdJeAjXm6azdksAt24QHMZGMHeBFCv72onko
7N+bf4HOY73bJ8hqfsPTHajGFUVzzAhCZRqZlze4K5qRVwVfyMO5bK3NyCxQjJsCaojM/EeiHKiT
RSoM2I7c2sWgFhayUps+Z6bNWX8/UQ+DJ+NR+RmEqOkx7qK1joqFMuRWAu7J1wdbOqma5+H/i3dQ
qP/3rDad+7gn5FwgyJmtKLxU1fbWN2njhGhat94OBDZs9mCMSZu2TnVL3kMCip6OzCFj30ank9jx
Xk/PVN+Is4AQGc9x1yIHVWdYXnvgqugJEVa/B195pmnH/Xr9jGpmdHTtX46fl9r0xXNGj5kGqqQo
X2q8rpgOJvt7yk9xVWL37btFjyS6W9mfMYNa1PmjjlxnAFmZO2fHTLyHv9MRs4BQmL3P1uPwGhCz
2Ibj//Vc7ZG0irnBh1xW9DJDnqozhb4NnO1lqJuqC8Anj4y1reECvSJ8gMy8ljGQ3mjDcS4IsIxk
KvCC0k1niAnahzEJcr344wkQeFVvAQulpw2EAe79ttmr0OsQ83VDtgAJLvUvySNtcCyrhhCGGOfU
R/LQ6Su6ru3d5hCczE8w+zvz8pmA/ZYQBKA+b627dD7Hyh9fC+KbdMzz3/3uKQSz1HNYtc7CFmM8
l5cSQwwaeMqi/DVtfXSGuWLbB5wX465QFfoGuuxMRPa9VT1v3IbkPfztvzDRpaVBw7qxmgYMKJ2A
Z/NPvxNf6OvAPfoDoVdM1YKjhUqIInyl9WiuQYfzxcZ+ULotfe8kGwCEExK/lFU8OmGci5Dz8B3p
AVpSvYChOPxZhjjiDNnMr0mdm+EJCiXevLJ5fWek36YWjp2XWK90qrAV36YlmNwflV40+gCdapvo
kb90tUkJ7V7qWMJ6I5f2CAmQeKp9tvFhR4uElLbHMNz1+de+R/uRH52k3ZDZqc4bJpRWQx1+wKLY
OnNtPo10eSHeDHFg7bSaCH5RPpya53PQ1o96siyhFL808eWUGPramWEcxFJomBKYBwBHNuxu3416
Ityc9i0xHk12QlGLPt3GGHXNhvMURGDQQhP3dev13WnDd/CguGmu3Z4WqEn+y7Umd8VqcUe0mlTC
Y1XVi6/epjc96OKgIYqiH9QG+pN1BK5ybE0qKPlv/qkmOww4V5qMJY/DS7FeYqqLpy6vgECeSlro
iD8MZzsRT3crp+fHU98ue7UA5CuoVipx8lG1s6LKlYjPsCsIqzwPU5/B265NYafMVYUB2O7YlWHY
2bDQKPe6rNoHfj5ZTtd+JGJknohvW8aCTsSso8xuGxw39mDeDhooXNLdAcagbbdvVSJ8A3I36tD/
a+MFNNFkEflhpu2LlmyO4hL9WlEafnCnQAXW9OeaDWOH26t76Q8fWUbd8XOnxvFxQm6kULlEpoYL
GtAT8BSVM2Ful3+YtOSahHeO1oRwhutySLux7jMralxHBspffsz5i7R8s0sbsvgqGQxyM3+QlJBJ
e4nBv83dd/1Gb3bjLBTm3fERjgcMk309Gnw3iWcL7dyUoXtKaye+PC+zsXvLxtsyfZVtFKpZa09E
XTMWiulXC7gO6EV/KdaN9BmySKlpvDUOZsbMYyEZkwsOws2WAdVZ3baZ4vFUwpJUcLaEJY+Kll6N
aHia2IJ05N4hSjr7QD4FMBi1PrQBmol88+IifuWKkVg2NbABMk4ruoXjtyMRF3RLO0FdKCiB+RIb
nC9o6zAiP6dvsW3TIkgj4U4shriItXkpbYDTQ+iuNoFh2Gf0FWS1+ksa6BdW0iMBtz2TaLfYvssP
ak7CF6dd9NizE5BKzgpqEIImocWm6qQyY65aViFVMJSprnxIxf52evh1/49mYeBDDcq/PrBqnjVV
H7zQVufnqWCGb/PNYIXHuiedgVEYRack9v+g9uth8exUPoPg5xPuZFz2IM3QtGjEppjcNaZYtUmV
ADKNipX/AwYfd8gRlN9BJr4VE3pAO9Zpz0z9H721F9dU85JjTk1sZk0PRLoubEZMpOhViytgrs78
nt1MmGhfsUSdUBiUhR19GdEP1CQlGhXs3IzBTq0uQwl6iZj2LHvLfj2hnKH2/k73rW4vofy3P4jy
JXvVnxHjtwoSrpyufGeXFS7L+acmaKGJ7eum1J3QY58trq8j1ZjqQliJn8K/wSLNcqEdkPgd8zP6
2Moav0FQ+7hdEmX8ddZ1nd9e1WfUfoay1xhr9sHBgMOeE8nBg6YL7mXPY8x4TVWPxMr2haVY4VNs
+H0L5CXuUvf48VscpUl8p4Fq31Wt7dQIXlbYfWwVaVSe4So7U0a3lcqzxfjjp2LyWQWTOpQfq/vE
XwbG5ZE7N5VODMUDMQa/gGOD+NLTmJB49wgmyjuJAcHR6PhrMvSSe5X6mKmpSiVQb55PmnKS9LLD
dTb/+CahGQlJcjq5eb1+BIl1Eded9TgwHUNXj2ZupQDARO9UhOtZs1YgBuxE4m6zf/G0iBJaGnKj
MBLe9S8gCxVQsIEVmG6y1ebdiM0AgNV7F8kjIki+ILnQmw1lwTTmESWR7RvDfdjdmMS8M7/nqIge
Ng4xhtv24ND7K7Sss2wdQkVL6gZFXh+mYlSBWbD69rQ/VYWvEbedAQjfbHcpB+CLC4ASD9smRrAj
dkDrOGO+EJMYjER2z8ecaeTiOZ87XocPXM4EqSGcWdWJrKt8LSoz75SvjpM4BP2rOWopQ4ftV+H3
zxx/sDf+UxxQhmMBLvXXExurxxxYO2+1+rwhJbr63qT73gmVxCk74Uc6ADcIk707MdzP7KiJeFb9
LgiU4TAgHBEu2F9TjghU6mMVvsIkQC8SQGbGxQMfGIHSfFixWJk5O0ym5424UV7vnV1MSua1wahR
MWXnTk/edrM0/X7NLYUtvRIkIBvcSU+1Pwx/E+lnz+0OJ8ebx4fLuEKycLjIb0vo8hz/n6hViU3g
0TH8B2a0NZuBbmUIJMo7dd8j0qK+1dQ66Tqnsx2bTcrGHQVx7o7/0gmwQdf5PZk7AulJysykRg2P
Y8iALSw2HLLv/TKUOEagPkzmab0chzooW5E0Ag2B7z1avcClW/E2mjyIh0wp1k7o6rjAn5iFRwWG
JujzPJxQWlGrbh7SK5QkXal1i65zKmIccszvCZAX62E9JN6eMJnmHsTynrxYteNGrcgcAYhwzHIG
515d7orapy6VMdaqeNMnb7GNR3ST5ZYAXLzUpOFPLwC/jgs/bevjwvtyXbfLWN/GoTdiudkNFrDZ
y2KZLhcdY9ItzJlWodo+gFCAoQ4uYh4r+Gm56Pf/w2PmFF4ZzS+PxdBs1EnVrJAUF4Dw8pRETlxz
BFk751z8ffQh12tCKyFoaJBvV6viwAjrZLmDh4nbZoZV8FaKJ7nC5zjfn5MynwYtASbShVUDhSHB
Q/gxvbHoDpnoLi8Rfv/dS7UMhZohi52kyGfnf+6zngynXbv0SP7S1ndUycpbCpeRnsFFBmxehx9O
cZi0nHhGp05AE5mxUtjCJFXBPAiDjPON4NFMX7xoXA65o712ZK6cN5Rc/NeEpiXfE279rMNif/hd
vsyiUFi4D2dQsGt59X3353q29+7rjJlnLaLCUTDqjX+5nlTRl/fHOCOiLg/i1Xjv/82oweguwAUf
wIkMUeT9VHASyR9qhTgTIX1yQZR261kCTOHjQJNRsT+OYOijH4VyAjESZae8Oz9TE+t3P7VumqbQ
D3loU6ieHArCgLrn2WlSFu1zDAX/I/kNbGVSSkXxsorqgpKNV9zFWlodt6Lk7nBlzI/wlnpfvVsX
lCVqz4+t9FkvHKyUSEhTiMPLHqtmTDyEqa99hgynsfyGk6Rmto/TIdtfTOxbCg2d7GMourEsKmEs
bRLOeYeZN0dYjaRgRrCjw+i+ejQlQ4ME/x7iu665ecx3ScYNktDcPVkWChFKUKeVpfXHLq0lECLP
nIntqegQCDHm0GhfrD98TpJ4VNvaEBCzBOiYVajmfEglexJu0j8vWe5ncLLqDMNyaCvShkBQfKZ9
ljepbtEaospAumg8+onmOPjPgVu4SVjG2AJqTe3eevXwBGJkuGARphwd2kZDIDKeUq/xG77EGNaR
Yr7llERs9tiogFGs20irbY3IuPC8uKmqG/0v1FrkpHm+trsgevAdApK5dE4+T1i3N7uKxc5Wc2e5
g2klLT1DRLVpaEsgc8SGt9H5myjFx7UoXzwJzb2KGSkrtI0IrejTQ2N6zP9IDMrHW8GpHgfsxVE8
FJdax696cZHbBcWY7XDugVJRUs41t06zK6BU3HPn/g25Z8nfHInJA7WgHYAc58Y7erdLrbivqLiB
vkF/W0FjJpxZWtp0gPlFtl7E8hC7Sm1JXN9JrEJjjLiYgnmA3f5DRY2fMrYN1DBcAFVvodwDpj/O
jrAYhsHHg0ucvr5F5UrsR64p3on1QMTmPprfR4W92uOWndRzGonLD43HjeNYqJ5XEsRHGoJPl4/e
++vgKBBlK8b9YcLdlpdrt7NLay/qF7/dcm/+0SCeX079fAT9/lhmA5Hofg/darI5jJWvqwyrVGWJ
+ebBbyH7weqd2QuPxv8P35q7YGxgECKQxOznkjg1MQLBeCUhuruYfTDRmcaMSAUvDEOfLecsMbs7
IP+Je6fVk8N2jQuTJ1e2FMe1hlhrhnS786dtYSNJz2jWO44jv0VX56dE3mFAscn8LCe+BtYGB8rW
AXpgVsgbHE8I62aWgWmmQVtDdYhySE+X06dGM7hps9fJQIE+eEWA1b7670HCQW9+g6g1gZo9k3PU
OWnWCzUOxP58DlAMV3SpZmbEPNJKi6RnmY2EXlucEEMKvQL059otZg6VFHm1qfX7mKc+RzGH9wsE
OLvn6q4e8rS/lToRdCJmpiRuAg0EhTLeMlD2AH8uX7iuoOqxyn8f+plLIwIyqLl9+5mlqx8OU1M5
YTQ5WKLqDo7wjsMFNMn/U+lLmxj57SY2/nRCVyYlZ/6k2ZL52p0N1NmTlYBFN4Huic61k8mm8b7r
i/Ng3FoEAtTCtF4IISqIY4MB7jFAbNpPY34byHL3b4DUTuMoWPcYaWlpShpHEbAqKpS5WvnlVTKz
wnCOE2H6WW2fwrFiJvl90IUYeAsqzGRL/hrkvRjbAaMvwwCRz2DmSARtPmUQ1VCDNkBKa8QQ2fLK
FUItYp8r0fb4QRB/ePAhteH4cRR064ozTV0Nl/wtY/WWxHQdYmbFIEEUAh77C1YQKqv4TneeBWH+
6JiSeJnnfZaOgpJ0GIU97OohJxz2Ntx+J6PNZODfpdiZ/kqoToso4fsGhab4MMHieiSewYjHZaT6
HHfKN8cgczFBjN41BmfxtLDU5ctAOUsnSXjEc1lJwlGWR02mLWAOkpOrSCdelkSZKiDiutPJwMkI
t0GA17sBCOyQ6pJ38T0YsaAyPE6xqMS0ZonkViCo4GVc5yK+JyM4nzYjUskh4tnC6Xn/gh02eDnR
mMnTHEwQjp+zH2NJgtML96sr1C+pKGBgXMlXuc2xOsQ6pFXpj9IKX89J/nSAssm71iNc/b8sbvOQ
sS/R/7eQdxPRbaJ2YFBye2wFmoZxoc0NwyvHh0hq9olKDiuoUMyarI0dG2Rsh5ao3LnuIz4SDRTY
MROedA5uorMNeOwP4ksqF9t0BTRhNT/Rj7bsR0SEFvy2tLQ7tyb8IU4P0HPtso4ZviSM9z8vpY6I
lRKGRVfrccRN6LMmFqTAQytzYz+lBOM+5mWGKZlMHd225ESOtugAoA8FYRddSylEhX08YnbaflUG
NKs0IT2AWatL2paGKNJ57eNMLDqJ/3obssjBNm7JtsA09mzXJ8ojN/feyK7j+dVTtExTnrjmFTLH
Xq84PbY2jTe3Ii80xBQuFzn8Hznbw4A6DxiymUVw+budIiWWw0KD9OyUSjqDb+7kWZMqFZIvsK1A
k16uNLsdI37RXSSmnoYkiKniuhihlrysmufHbwVtsD34Oc3SvfzfIY3ldlWPuJuFbf4R9dJoQ07f
3+rwIz/sf+qBWQfMRb89WLi4v0bSzJ719htl+wr/8R/d/LPEs8guDRdhVwPFQhZh7+jVwY7oVhmC
mNdNHHJkIIo1n6z/88HfaSc/A9oQRbP7gblrl7YxR/Q9VHbzhMTuDGEpvZVCGS7Y89EXxjKNR4xI
vDqEqM+LdFn4QxtRp+g8IK9ZFI9TIvtMZYDzqhVQ8YIQ0IUVJlKbc4BMy26c3uVHxg7vC7NdShzF
lp9q/luRghGlJWCNisappJWErFZ0nR3SoOeDEDWaNTiAx6QFhZQ7NA6qPQb57Iy+bfp2MC9poJN4
jT3dwFzNGa3bwh//vWLAKI+pL7KE9lF4pIdofJdikRP0ipnGl5r3gdP5l5U+ZzM7636XFlQDtHOg
f3HTqU6z/Nh0IboG0rtsZP8rUk/843YnSm7CmF02w+G+4rDsded/6B6NbI4QB4VahpM3LgWGYyrv
6NT56Pd5omOZvVkynzURzdoMZaA+hsgml5nPyr0RSaG/5+wRvZsbpJqtTlDAKqy+U4UtRJNO/Qrb
paVFa9Qu+09ZQUuORroR7hLDYhyVI72y2DeEOuPjkV1PtIioITywrOuIwfC2JCYg4JvBDdPRa35D
Fpj1b5APnPy/sDcL1+NFsGobvcCvm8SwfhFPmlRpnsO64bmPl/zD2g1tyJf7aHS8PIAdLBUQsFpi
Jk43HLiWA+dO8BVmCrQeT611AeWXinhFzg8m+x8zoDK3Cj0ot8MKC1NV73Q5YzhTf5UqA5nAboMl
3QtjcaNXv1lakpsBthi0xmKi5ZBfs05JL5vWvAUlT5W11KVu621X7Y9tf0kXkGP4LOSm/ExEF8Zp
4xL8Kh5ezc2ZEM1t8e4ng+m08LBIVEMvdxBTKH7mrZ8VmG6aAW6R7fCKnpRpc3ZijpG8HFLETptf
Dn7UDBxe2v23mMPuSx0mOtQIwxYRladirON2NtCqwRt5KXvq7OcRyhai4GUki+oU1Dk3gyEAZewU
XQ6SDir7VnwnWZAh/F5uYuAZnFmLOnDkKAi9HKZC5S+qn0zOmJ2AzMCKYVdLG9we/dTpcUOnuU33
Wr8KZmKD4aMnoJQzRLv9yaE1q+hl/SUqS4P/bYu4dQ33IcjMkERibPgna6BXsPm3e+h5vRiF1qc5
MV0d1D/TqE3eDT2cZW+Gx5Hg6azQoEyKY9DsMePkb+9knB4cTMFSbXL9yuTjOjoBdEmvggGCw7j7
Z+ZZp5UOxhXbP8iTF1e32HsvJ82Pkhg/hssOVvFlidd1ucpmQSzeK/1jOLWSlugRhDG2vLboMN0p
Z8DWk47f4a7S1WL1S7JgsNn5rFOGGmo6tebF9oGGQWMq9vUtOnS1NaPBYxIcQGuNeb6hCgq2fOqN
pXhGD1jch/aJ/6Gjohj6hHEGRABnk9YeHt7L9BL4N/tU0z5pRIypohszRdhGPf/5b7plHQEPQ8H4
Q2ljJpJDkYdoj6lQvewmo8iXazRHR/+Sjv42RC0oU3jlZ31FZmsqqwylHrMVhhz2fJyG7Ik2zsSv
MmqFvLJCbB5KOd11/CUNNiV9EkBR+R/jTXPd57yXssYj4lHisvc1TsImA3yy2goC8bgPpWcnUexJ
G8pTRZpj9ytNRRdWqgZ3+G7Tro5epsCZbKsel4SUwp7wfCWKCrrL5H/08CcRFX8qf8gne+6lyq01
JqrTY2DQ/fvLuCphGEx9fX/lauBg/m7/g7xjRtiaAa9Nf+l7MLJv44rmeBZJnAYs3S2xI5BG5byN
Wm13/SRPEyXBMikgEqK0ID+aVFXoT06wTNb+qVpor6fqKK7QacOcqtoaM1w/vmoRkRymXk3MxIlF
lL1DKOZcn/VjnEK+C61HRpf0tOYJlIaXNH00N2xWJhfJGnPVLoJ1b5FmzAcXkgnJb95okjFoLqNG
4HdTvCRVU+ozAVmDF+dcOpBS+NDtzPNGxsHTP0pawWcRMD9m1Opv7DZdmptSw2tCbPf30ZLAdGU2
SHHq0Mihc7xxvxLdagmOgAtiiIgbVBpwvW6q20UPQAY5Xv8TzqK4KFziekavDEc+MbiNV46XcM7m
evdL0ijwaokhxubygHGF0RLFIPECOMyCLb7xQlTqfivTqSaD66+uGvcsovfQoghjlK1nuzXWKZx8
eGHaYNjHZWgZtLiHs7ketPxrbXOKPEsCcvIJpmINo/qmd8czaI4o02DJe5D+v3yG3gFRGPCC6Vz/
VhUgN/PDqNgi+JlVaQKHCLfK+2FWLcRJqyKq6Lpu2scfMTQhmKCf7kLi8ikHFe910jHkFtQ+D69G
wgZyA6G+Q4+ygdQLgnzukQshM8W4n6fVWTgnVFFgh5+2dsfr/NcWFBJv6Znhzxted1GKjHNAMEU9
WOYd6LpYZtGZAOA8paHJerz+lLr1p5kNwRxDEFp3YThUZPI2g6pvf3FE5Z6gQlyyPOP1eox1ml0X
YwLFqEkiHFZCp09xlcws7uYbXflNhMCB15hHkkMYzhEoPfzNFVWWLL72UpyWhrJ9Do3HrqdCmF05
sS9WYaE+IeT7JDEskMOGfJ7z1xTiTQo1PAuM4JC+G/Dc44cJNJPIHHwrGfYpQNAsXDh/My9IuWbu
2gkuerKzRu1dwYTlesACr/On353OxcqL9fDLlmJ6U7i+hDpalNDOWDVM1LpWeeg5MDhZstEeTP2P
fsQvc2Pmm4FlIPS6kYBVL1vhUzdjPs5ENJipxBR19yIciHAjmM2vuidwGQWz1SAqppstaBPnGrOT
LJ060d3iD3DCxNTTOUbGFmn8S8u1mrv6XksCcF78m2SoBUZdNKCNvyXyk6RtXs0rH0F/LJI/t6xd
NBUnFRtOCNE6/hHPakQTFXEfsz0UaZo33KypjQmyQvf+xnCgz+kH5b7Q8cZem1Dr6+DDYbS9ba2F
1tyv3fb4XAv6fI1zV+wpqQcsjfq/a2et8u6sOr6tBH0IJZzB5CeUTbmf2WzLarV39RbNDrPa3wcn
jXzXu7p9gYN6LTlJ7KI/lgAkTEVaS0wzDlaKHjB/3MX69H1G1Rs0NPgu8XHpmkWzEnhfsBBs0B+Q
bB1B2Vz31n3Z/b/E4a2kWCvqx+KQTVFTqLOxajTvt46mkQNOi/lBqyV9VuNJf+WBcmhidN7fV8gP
u8WmujPJbuQ/N5pPKZRkavBFKY8IrT5Ceg3a3DalqiVnNOOGAcsXtkvl8D3todYQSfPwB0rCTHEc
2otK+q5UOH9NEdaOz98MiuiZu3+EhoQxCjHXB3cAsEx35BTi7LIBRQlLRktiN34LR0ah1I+9EXo8
qyNck1nzjpghWSuQubg73PrqjXEFq/q4h3YkkWLlcsH4OckSGGYEh0uxoAewstl4ruHErra+9/hR
nrixi/uH58K7u1I0VbehlnORiulVDyU93agLc3ujsNQg/AL9G8gXqq4fbuaKgMlaB8Um45rq3pOI
1qAAl1oc8yHqsPUze24HasoZr4tv1s9nzlyKtLfnnnTW+Tk3V+f0DDzDzODIu3WGbnjmmJI/wDyM
Go2tpzqR+gMZ+L8ka/+rU9C1BRdydz/LXniH2fL/QpbLBiDDHbF2jquS8xu2NXOqSC4uES8QXlea
dPXCxAApTF6pX8XpqqH986Wl+QT33nyUL18Xv/8HixN8RHqjPWsql3+HLPnzlJRgtFA/uawJ9HtX
VOuJ9Dn8uFkF7LCQtpMUKCgs+oAyVJKxandO7KmWhOebmeQ42ktrkSLiOm5uiLkIoM5LnrgJIHW4
B9InFQnJWwWvQdIgvh9QjXmxfUD4kg58dZmejtTmD/JTU5XpjIzRlNIIojGvUfioZa2I7H/SI0lw
msw4YWzCxstCcW6OVECaB9Rn889PBBLSaCqf9PQe6AunChAvLy20klmqYZqIZau2V1/c5sf9ZnxU
WjfSK7EyutcP45E604K15U3r06B3BaWq2UnHfDx/uadcvhzTL3qu6a8dr8R9W5tvmSRJu8W97okJ
lomNSWujoo1k/OOI1wVTbXII49ZvPVu1Qgh0BYXGb78zpIyX83LtEzjFBQsUgBhYK5/PO81FV7X/
fCh1ciuR5CVNcHDZ1en6U1jlhfRZRNu2kEiYrtDRm+f0J1icr+r5wWrBpou/TMnXolZRdTnPxyVZ
Zk2kNkaKRos2jJbSodSMjaGyCtcuyD/UnCb5wUy8JgVzi2rNZ1r9Y9Rtg11nHcvX3hAtIPceyiZZ
vgPHxpiIGiLGwlznhYawl3Mwx+eqsp7GYh1LV8OBqWbj6tUPPTH9zFglWN5MIoBXXG1yO3vkqVM3
PNp/rLqCy9HnHCkv+kUzH6vZomGJcw2eT0C0Nu7xt4Vsd3DV2rISx8oIEaYxBpWvsC4ES5rkaotC
ueMDCWPVnpd/C7OHQ8yI/ay7cykEfSauOxJM/Z2BYHElp9R7mKpBWlQZD/nWqwfgllFtn37dVsUg
GvTioAgAhhMjaAAJLit2pMBJWdpuclbnmX5fbOXsCMFr8msgOkEtSha/XnCc+v6p+8/FM9zxc9nr
OkUmCHnR0lFloT36GM7ndxrLCSRbm+cNZyfl/QsYaH+4J82l552SVos6jQ6hlOOyihNqSeW0NvFg
LkXFyjVPE7dpXbkxRZHQHTBD7/o4shW553GBcmN8v8nMYCRQC/RrNixwuFIoVwDYXvgHa5g+s/2h
hEcqFHoMvi5ufrccP7YlJiYDCUYMcgeOg8AhuQc1UJBX5usrp4hdCrK5W/wnXgJbQ3RIACqDwo3S
qcS7vGEJmfPzQLQ7B1yz/y0h+HUKYT8NlGp/oC064VfALxv0F2Zx5ROzaUkjvuVUQEdkrf8kAzkJ
FSV+8VzLkTsK19a75qfDCZlHvDcrmkV9u9K4scOv6xmZ9ZdQ55A3a9zcpYKKhHj9SNs0v8pMjjdP
Za4LEyBdn0xl8NKzPn+/IhtLEbNAuOSvd4Y/4WWRuuxEP6JARkDciuv8jWsbGL7SSqd6CE1jaFwo
e+YDtxT+oK5J+bZ0wJTcH8hmjAWHJ6jPXkrqvvAfMIpAC+q+LOOMdBAEvwja++kK4QZo6jt36zzp
Dd/ms/w7+Ax3jte4ODtAzQBCW6qpFnIRZxoDHVWjhl5iIK6imtaJ5zkuuQfX/9nuIG3D4fGPlwan
rUykUnc+0Ou+uoX7xsI3blQr0CgpiZe3nA4cYBN2HxWdUwAx6DsgR/3G/hNd8e56+L7zVLEWueE6
njYc1S5/i6YXsQ7wktxjGjwaFZ5kksvzTTUXfWL3INVF5UVjbHTIAmDDolPR6v2VC0fhPBJp4jdE
/teg1I1ffotAZY6kSmJSGj95ZI+1mB8+hpcNWJ8oB39DK1wPIf+bVJSX8wpwmSSeo6tSLVZeMxLg
OFKXpADE+iiMqex/W8JyCYhZXbxjmhJ9y0/5D8tmtiIGVopPKeJch1Qc/HG6obSvroT4wocVpymF
Gi8C01iMBN+xowJ8ruDom9L53RFHf10OIs9ww38dqHCt4y2gaiTtiRqfqAcpI5veaZSeJNOJZ22H
Az6iP9d/NczUkVl/MaxARCoP4qP4GkCG1m9WzT2Au5wTAOxfxB2NYmaoZzafZP/Px4LYFcfCZ6JN
ku31oX+NVak4jEO6++sJoRfr45vQm629F2l/JwS+q3VZg+2w57iB9iQXk8HLRocD7GtaDwRJwhb5
RklZH2t0X/YuIB2u+ubdNaS36CuffazOVkUOgBi9fXcsKIxod5uO/oF2y3rd+g9e3KBmMFiZ+8Xq
NYaJByl1y7uGu3qFEMVZxRYCthyUmaLWDJ20CcO9mIBo+5/l901egMi02zhWZeH9PYRZ1JaQuucw
sEMS9LGbBaAiy1ZOns8ctQWCYIF1I0jLVGhTV41f9Q3ANTo1GrhKKi9wdqF1Q667pBxWiCLuzEQ9
Rv3+1RGNoJgTTLUw90R9MZrcRwTUSdRB+hj1LTnXsvCjh3b7eGPhXNpaGtDPRpsoV25oFinoBVIR
t67ZFTOH7SSoaWIiq93jFsreaH/GlMaWDDivVrPNJOnQ3eGVS2qVVnMUr5eepXuPOTYNQ0xUVitX
D8WKP4MwYv1QrUETiIRR4Qq+pzqw4aqH8Pkad8Ei+OUiJ8mGN8S+C/dhKOylDM9LeZB/zabB89q/
x+ovKbjPO0P6wSzmoMXSi4aipE3sSeJTDEEKCsXS1XF9ixUaUKjurXFTSWX7c+QM325GRY/p0c4t
kecDr3IbhymQEvXGQobv6dYXdxAQ63/cmTl+DTk42dAiSN5JCTAxFD+e6Roywg6bkviQOj4k+PAd
oXl/xd2YPJ6onReWv1rFdYUnlx9SrR2b4mnNkJbGDkUOvpcD/cfQjWrLrwK6BoZf8K6uCLuUoxSO
SKiQoqAC9hSsvq7vd8TKFORTdTePDWLD28pv4+5DM187a2z5Ri04yjO9jHajEmphFYsg3m+Em0NB
GZTsbtJJFn6TWg2WkZNg23iK9mTcXQwysnG6uAlikUdD6QGRqBSjkPlRFmGDu4jv96G6r1P6TVnK
BIlipcVzw5rtbgeYdptCQod4jlpmTSBkswmGZ8bXckEh8BVQMZiJ1v4Z4pneNAgw8xAqDwZ4gsHK
1m2dNAgXpskDUAhIoty/vJrjAC5UI4Bg/S9iXKgiCD8gkGCW6k9CJGGY9UErlaHhwntokCgV4raz
BfrKImIy5nJ2yAT8FpoVHJEHvsrwT7C/ZAILYB/hGZrz7ryV1W3qqS9tlg731OiX6GJYqBgHmepo
aeqawIdXHBF0OJLp0apLLuqQBYVH/uLnIwApW0Uqv55UosoLeCkk15HsJ5OEQU8Tn7RP0OwzaG6Y
Z0RatkdMF0jWNl6WwRcfaxUZcsYmazkXGDQD7WgHNQdRf/ULMKq73+AUSf7tepNW7OGiiGYLWLoR
GAWqhkBksohRVSSCMx06yR3yKF4TYha1Ty3voQbeNO0XdufdqlqjtnYtG0iwPuv+cZVClfzBakOp
7gQD4wQC/Y9+WbmNpnXlF3oaQxqi5QdFrx77SE5Dw0UOwp1k6bVhX+kJPHwvY0UhIFsrom/cuuux
7P8iIW59LzrbV1mGqQucgHH9Ops4xrxcGSl3O2NuVzog8qSQiV7QXvuD9ALU7xpR16AMuxa4Pbns
8ox+hw+a6NlmlSQJC9g6wI9Tl63QH/xhFFMTHCO8Ti9mKvJexdrdxIayfVCPsV3QHLLP7BC1wZ0Y
qeOViusCbbgwjqHMhJIg2MibU4diCwRDlB1qvgoZx3Jw31j9ELaVU4OxrxpZzUllgq9xRw/qFete
04P2dcl18hnxi69IvMy7usc5x5c6izoBHlc8Y8R3ZcMjSAkh27Yzufpnn7G8RdX9qdseYe8vps5k
mAsNTm6N5lvLD6cOgyUuT+TbUFBQRYkwAJNURgwlVyEBgeNWxT5kFKdZ5r+IDkGSq42ZsFn/62VZ
+bqozYPrcNos+p/m7cmGIeGMcw1L+o8Mk6gXa4GCfFIkeZg+J59TrpBYT1R0re0QP2dH6v2SXm9i
qeHN6jCPj2dH754WMyZ+E61V5OHB5mxbj/K+sfFQjOqDGTfNG9KAFJDq9Yw+cH74I1JYqsWSmURC
TbWUJu7plT/+JciDrXqVzZyHe8BSOOVlzAfjcbdQ9cAFfwuoN5UHXyQe1D/cbXjKIYddpyw983R8
NK68tIFG9AIlzKd06C9QDE6ZwOh0hmVP2c9FOukIrzZyTp/GE86GzDYecQwjv360XlpVd84NaXt5
u7IoxHVVkW0A15nfRVc1L2NSec0lcPkyjnLX9okTWfVKhKDegVc746dGf5BPWwKYCRGwbOm/FX4n
+yyl9AW0Nf2vTxhZLCBnn9rz5d793w6Lv5XLvwvCuTkWl+cdVoy+Rw5LHNFZcKgJCBumMPqr5l97
jD5N6/6n0yU5A0eqDrpokHcQvLA2app1sYLP9laysmTVdy9cUJs0eBh+MwG3D8JlYi642c5daheg
iEqKEQ4Zb1KecMQlxtnSqgWKfrFZy5KVOSq9EgHddy0ljRmPe9fTe9JCRlS7cb6i0iU6wx5IY+ar
wrUOrH1+YsZzpt2leyJIWgEW11Vm/WJPMJo5WEAJ1lBDIoRR5u8xmlz3cqgTX4NlejNBAGD0TqqU
1Ivpz7Tsy9u2i4pAgboSzg+OvgOg8r59ecw1VI5qodce5JYKa5BBs8vulHm3EmdaOe9z+LZLxVCO
a1UNF0V+oNl0ftj6ld4VEuEnAgBVZoHej6HdLAZiuapmMtZyJDzhvbncn/XBBMBD6qziHUOn90hu
zMmD5bQJzpBBI5K+rNN+6Halw22oRJXc4pw6LVZEyiQFOKvI0UfMkdUEF5t6Waj8FhXM0eV39Vb4
1oAjGmcGSulyD7bLD1Yi3n0x3nBcFvQjb7353iV2SsPZ3HUZCvDIwuQjIxHhY9xYUEM4ohcw0KJa
UxVMGKi/dSWJH4SiXfk+0YKkhmoAm56tOrnrEXmeY3KxzbB+3ga7jvgYHM9rQgR+S0QYysbtHxNT
861JdpxHfRy6B1eMkTpPM54uH0KESQ/ybnKKBQnFJepDEF1u6Mr9AS8Rija1x7DwN9MXAroffdIL
x2wgachZ7XwLPWBY2RhH4OFzEmrRJs2ZGesbB6K7LWIR8IPBasV2xpebnAx7ph423aM4Rnf0yptm
xNbGWb2BOD6STAvrY3wY96/89EP1AkgdIaBCLTqsKGPMeU1i/hWvfC2WuEaIZdY4a1PTNBC7oyjT
TrZj2JqZBlhxgs6wUGchwylQ5v2YFREPyvbmWAnJpjXpSdI98ho7UEGDQMIOCvpGkHLg+2v+82nn
/q4z1eVipoZkQJOMq1pzbv2hTNLO1L6gPXnKU200MnbuS16KH3A6qkpDuDcA0SDook3ZHkwCTYvB
0kOAp6OHTrMf6OocZXc/ZQe91siZUoFYK3XrII3W+Qkw+OA9oJsDxnphclH8mhUv3rQ6w20SVTGZ
DOs//XTwcq02Y8I15Hx6ynAQfUp4wCfaJCetubPeyxIVyfHotQUiufmdVIWpiG2U3uw4ZG3dTc14
GvSqRS2AvvPYWS+itydHOnZtNazRMB8gYnmGZIr9hwQUGHf0Ap3DmoFMK3pn4glvzumOUMkzTJ1v
PsMcve2rgxGXvnJ09S0vJD9aXEp1iY3k8xo9pIckfhdUtrWDOIv8S3jFHp/35soTrB8IaZDIch1Q
fD6ypMDC4P7nKh5J6RhDgUBYtryWQOEAmvXJSYnX4EfzRlqiIFk3N5y4q8kZxmM4AyVwG+vr4Lji
RsMbfPyQrIpHsQDs/JLeE0JSe05+z5KDvn6hg9Kgu32vKzKyZ9oedQJ2qtJusdhF/Ew//fOQA2lZ
b63IOgN3dHqw14d8v1tkg3ihL/7ZTexyHMlLxpHnozb8MPtwoBPyzr6p6a6CX0Syim4J/BPH/oZQ
nIAKz1R8Qd3AZmBtOIYju7gQOGE2PlDyJmGzTuTjpoTK9S42ZYjINrAkEW7gV3XnHUrpleeSPNzn
u7U1Z3Nd4CbPKy/TrwujcIu9BNGZDUhXSQO1egpfsr2EeQYmbOZvk5qGktZ35uhBrfx4v5h6/ERH
VGqQjzkb97wVF9MwmZaG6bV5uT/g/aj7HzMqueC/4mrd1Y0RAyCio26hoSA/Sg0IEY7yR7HYfgEQ
UuaoHCa2Uj4bn/91t0c+EoBgK7JsYCoV9aevbgQ6E7Lk23rEgeOdrBOa9P9ynzXMJVBrZ8Q7MmE7
0Wr4Yc2hNE+UES9E4Zxg6eIw2FLou0NM5CQ81vBlPktsvzw0DvZRtwa6oM5ALAf09pry2xcSUb4z
uEt8qdBZr0gaNFc2jYUR9ejATRlXuI2spIbhP2LWVGhIy1pnhqWJEwse04mrRVAo+DuP26dEVHw0
X1cxCBS85LbBcTxvysa+08flv17P7YdV1eeSWL6NiG++qBSnlgbYsXK9uDAfJiK0tO2uMgyFylXz
F+jmLXNgcoLUSAERUB+tmvrOXzuURiQFCHruf58pAt/CEdVd/VXfsFXf9eV+SbH5Zw5ZwBWOogGQ
Mpvorm5gqFTaPcUGwRaUwZiRFqxaS0dcsj3Vtga2zpuA+J4tLj4aNTXKxfhKRLqelUrvhAKTC11D
s3WTLHg5Vn1WxGbWkXckl9fCUyAuXt9auWT1gAWSj/99x5wqb28kxYA6MbM9ohZO3/ixx/avuy4p
z9hCdanQsE98yMDahncAPm4bWvQfFvPOQ/iKjsEJIpXoCJFpCzyHQ9W+04HW8HqU+ccPBJ5PDWfm
5JAzGPGjcHvSM7g3jVhFXUUZGs0fELmWsqoN+XAckldl3ekxXf3cKEJUgMv9hzStyy3mZ06XoAYl
DGwjE59dKOWVj0d+F/ZF50xv1bCpH+1KxtHRqcuG+hsJThhXwosvW/O14cI/K7303DeGOyVZGP8Y
Jq/sgagQsqF8gjDURyp//5yxH5S2RyvBs6kXdPVWprY8VgVSxmOsjC3pkKDrGMJ+p/ubdBHRY1cK
qmHrxlxtcIwuYKblHVtJNgwxixgfVkgp0BodEQSwl/tMhVTS8te+28dOCHV16rG7+tKvJI5dXptF
KzYjRn6z8S01rTjwFRADcyoVtLQdzTjtrPZfLOHifMnYazLwfiWUslVQIaSBZORu0K0k26pLikaP
/sG8YcWS7Z7O7LK3Ky/WOA6i6X7Fb7xllnGgCYON9qWIqUgFdnLbRYRd1WHEc3l0viBR6opqQwrf
vvZvSoU9EqpSgX+NkWdBD5TmOU2Eu1OrokYj5qTY3wTldbuvM842YkkCZhZZqq5z14TcFwo5tWOc
3BO8O9DI4VdIexXm1MTpfEZEwu+ZAusXQfnKRrYm1RId2MSw/gH1oeBGpdV/3+zlJI/mRi6KEkro
d09OHi36v67mnKefqJwAngDCdNUQcK4zZ+gbhXVrUW3rU7iN8fKSuUq7ZKfR3TS9mqKp0t7IGrD9
LU3f71k23y8Uwy1q7/lFdOMGERIC7TLldYu4yhFwLWRV6ihfp/TDWjPkJoek7sjnZ/DOVG7sGkzI
sj/09rEewXYomcR4n1GoVFu9Ijq/W8dFUneWsGQBZ1mrP0jCXsvC20O/kEhmtlL0oZqH5v3FdYYA
YFgL87H5uoyrMZSJPysSsATDnJMwFIuC0w5J2UKmsi1NS3td9nfmDqVATVia8s44HbZv5uGfYFaZ
gn21pW5bHtfca60NXAwM9ChqT4v0dY43VTEO9Xd9cKANlleZfpcm9K5yyIfS4KhWDRj+3vWbQO9d
/WGfDz1eDe+FKCsW3iME/b8fpqQzeS3QmUb1MoVMj9ZtpsL79mFjlQRxsjp1/qjoFd7yFOVJbuNs
pinHO62SYNIwRgPlr89tPnDBguIUyWH2bAtmSv4MuT8Z6OiKg4kxrBv3z8kC0/tj8gGMU2B4fGaq
DLPl7WZZ/vzBwZ/xONmwll7/VYa8NHImcmMMDYh5Ygoad/1q9phQCkjNYHhtVNVWPuxlXB1nKcZf
nQEgddkGVvlDdT+P8gsI3OTLD0N4BFM2ObKsXKs+u5pZG2z2gx8tiknnkocc9qFn9Ucsg7pdoqqL
AMJe7ya9KvYlssWsebpzfhDV1dAKCoiCylkLsHqkGc+inO1/GQNavbHY1K0paYsVfhXiY2As1oZG
II7n9shmp/WsT0l9Hz0W7Xxg/2KgX1b6DQS3XgqyB9Q393kFsxd06ptXhYQwfybAO71OAiCQSPma
S9/ogwurcQQiBKrieVcu9sXwed3+O40LDBnhtgJAKAJtVYQqIqjkaI7ZsZHbFg9oIMO+b/Fc45PX
o9d6lpXl7EX8k9I1hiQ79BT/b97XnHQ/JXdoZHO+CPDDAKo269aSsEgKsGvNOM8HnZLy92iAEthq
ZypnqU3jHXR8WNPcCk8xWBR6+DM5WScUk+oQPNpnMzdf6f9FohrvNjruZg7xjotC0HEJONhQXaNG
rqtLxlEuw4BuVLfOXi1Ir+oF/yoWMroybtJ+o99nWm/EYvPlgjAsKTajaQgw1TKYb3SYUqGTt1XU
UyTqANYxjtdIg13pJWKhs0EjoBgH2jIvccQUdFIw4p9hFbZJsFDO+weEP5BheAirANzvUwNa+8Im
6BRMb8lKX5jTKEZIIdg25dPplUJkkWT5ZR2Ycb687jiu7qX2YweySfv9oRKfyGXqC8IYBRKX7gnO
z8NXWoO9fckmU+ecpU6BoUa1auU3XaRmwSNVWjawIMd/oO7QM9I1VSh1kYE80gzOqagAyfLV+NuP
m7D0gLViNM7aKu0cBbhfDfTum8v0IWW+SGV2/PwNPA+SIFyA/u/PTOk6P69gakXDjWQXzDcuV04j
xZWd3GmYDdAHLf8aJXM9vkT2kaddFUNHewjAQAS4hZR0N5ECXR60um3DC0JkrVkpniQQSxbnY0nS
KsAqx85Hy9gINJyp5HX5A+SNxT8mETQa8o8QgnQDVhloMjw7FA3jDANrwiXHxQb1EpKI7/f56yTr
gGAoKa8aUhfTwWV2ulwvrpI6fwSKhycWDg0G6HBSRmlBuLg9Q7KLhVqzu807tWsYevBaO2HGaVmz
iS5bRwbDGW2na7N2pZ9lAkosyajmKezhDmz0XeaUPJRyt1APVHTECEpWGZmqyaByao4VrMCgognn
V+quzmwJc5gfboGEgpP/TnhdtCHoHjUhNWR80PdYs/xOXkYrLXJs3yRVFJRlX1DK6x1JSYdaxcKg
mDf5fCxDxtE/MZdtiz5lxnr/RtIggmc4xpNYwi+MaV42yeLH2K1zxTQqPbrmdmSpry0Xh9VXwNBZ
0deo7N8DIP3itipJjaVGYHAhYTs4kLwYQgaLmYf88dGLh1N2LWS7yGrH7++zenQB+kqXIr4aiBcV
/Vu852/wBYvpb06MAC+VR0wqEEldYNegIqc8+ThNYkANgYruAJ8OsUq6I6sQklgG1B/LWYp8/+BI
4nKa4CqpWZ4chKdhSTLcsS5GGILPBq0Bj/kyPiILAiya+cg9MVMGRDWtOVsWUDXqNnnV/lU7ew9l
58mGwySVnmMhnNmd2qnqqljxgRF03Hdj0eLugAA1y3h8UuBq3T5RIpLVKXg9YdWBFpHG+vpoAR2z
cpaqxVRyUAbmmO+/z7UP9d7KULm2Tskgtxds4xZ4U/jj3jaW2hDRUdQPwrwdF0TC+Lq5DX43Wgxu
3mOG4qa6d+Oz21lmz2bfHdNlJW2xNj5r4SZj7T566/tI42ZLNTxHL6vQtsCDXczOpJhvUN2Py0fk
HMsTWaAo0VSh7NFqy6fL0za5PSq2PMpJwbWkg5g8XdHMOlv2IeVg1mwZg4h4utLgQs3boVNSmClB
Zkdc9dhoVrGgNCZyroapd7/edLh9PIH4m7LHIEsIBP4WBcJeAjQAttu99xGXrgOqDSH2R2E7BJl5
Ie2II7HhPtkTw1xKYLVVRK4LcE5jvtdz+uhIGXF0FbdBQLDao9TRaAEFcm/TGx7fxcS4sdtr0I7d
dZF6HDmzVUUOBVcOln5WNwLuGBWuznIV1Ro68hRHvH5HS69u3nLz11jd2OwNBMIvSSkCtfXj+0uY
cuBwJsPXP8ppqa1p669RSxWjyOQSn8SXVvaWZpyQzhmsNzb+HibW9dR36G+yaqHXx46y1Q0F5R6H
NpTsfk2THWSCrxwf/xoWqv3qZ48UqHX519mr5EmSH0cbnZhbxJNo4vSOua48MqBUGRpZgg9UZmqR
OAytdm6GFiONHARHOE6vO/h/JAnyU28e2pXERposumVfFOGUp9oOGvaSys55+lak1MdTtv0Rx5vs
jPlKJmZGAHxpXHUc2K7w1FMNzUlPvPivUfhmzsGXsuNxkfLE8EXuVb21OfMf8vuEaX9v3p0v2S3Q
ZvlUTEHkd5wBooI73C+fLn9aAmdspu7N/HI0sxT1cCnZs3NoJIyW7PMhQDmjB7GPVXp0SeTlZlAL
g8lFnGLfRyDZC3cQSLvRy7d7gAmB9Z0OeHoVuQniNqvSwuIdSZOvza9VugdNF3QY6KOOoX5idlXr
AV39jDKPcHKsewLW3dr4ooSLUInBJxMKE9zDQG33L9D7GgacCO5njwOdAyjOfuHKIZihfGn66iMJ
XYmPVe6ij2qUYRVot9uvUj/aj7D1iZ++Pll2mlU7vziQuw/ERf3Y8xdguT+hp3pcoXq7QL1DePN0
+AzbtTJ6vEnxST1l1u+Dt9nbwiNNy/2ESYGrWaLLt+nu9FTWWg/RK3SEmsRJoUhbgPCB8m45T3bi
ll0zS0CRswIARAnVrDFM6MMg9YaeNPLakF/v4Q28A3QZ5KyG5UslPi3BZ30ot7tmUv8O9eOzhs6K
he+DLFujUcXsVHMvjS6zCD8Vg3P51BltjWGs3M9fF42AvOQAvGFaftq0hklcfZvp4wseYUnzNTcg
NDyI0vs+GwDOtTffWEx8s5v1/rmIUE43yjl1B1XWCx4fmJ/qrgUAlMywdHRIbcdbAd8nI2TCvvHH
uFfiiFR3pLTbukjNGs0yEkJc9ofJ+3AbC/yjJHTkycAb12Q4Ehpfsa+92H7V6DeEvhbauGZ0TJ/E
Irvmaa6zFWU+yasnl4XIJgBa4qY6vpKymNz2lkT7j6qFQKYYXXY/HCnGlk0I1ofJ6anAIppUbT1Q
HvEpr+sZbySuQjVYnL1ABifj65KixRSrqFq32zwJ62y6EZTUQuQIrL+/mgqjVix/2UFpxBoRoENP
xOeDug4Mt0lLGcqh8H12a51KFHvYaFGRj91PKtXk/2GW1nAfA0rvCfLmY2djRwqZBM/K/aI1syCO
wNrhn6vN3ekKGhnVDY3msjGYq+AQN3vitDQU1szZX0xTb8MjzOXX+ZmRw4+HbjVAbGwJRftnq/9B
MLfIF4dITWj/A/dSDMovjG6NkKnrJCxGt+STnG5NPQU+NqtGTTNrAdcLdH9DT3uSL5l2QKaWDkqP
rvZ/kUpgfNhBdUKmRfdm58BD/3k8tYJsTVzAYbGfLaIxnRXib83ysWVSkYtl/Gu/ZUxIJzrhrgdK
MoxUlI9/dxONpWa5cATgXnxWTeNRRj+CmvfQxFHLDf9TFZLs1n+EbP7RhG4MgvvpWoXjg8fj6rTW
y8kFiemsLda1q4D5N7RMJIRYnaPPexlVguUZ1FX4pKyzwpxde4+A2vKPhi+gnsEnUaJ9j2KcGiVN
uQKcQCAeGVOuSsIRTloyNDmkbJHIlOd8LdzUsOV+1/ttbuRfhFESxk/vcevHd7/9ReNKOztKBpCm
VpVtZ3SWn84zJVQOuuwiKzFeA6DNBKW/z4J04qEuSlHwV6aVNBmLk0RnlPCmszEDhGTuGg9aXoEq
mwag6ySZwiJVir0Zb2ZwpARKxXg5M5GK2bfz8NtQVmtDlMjf2u7CXzVeMw9VK81Rl8d+oRX2Q34T
lW6rUS4dEUn8kOaVpJiMF9u/Vus3NUsCdKhzeW4+ncmaq/1gs08HowsQbbxWGYORuPRslbEpf9ph
RPzz11oLwULyrsSB32qLsEn4GAPUUag8jT+mgeqPKT3DcpCSAlm3YgsaNntoTWPJuZzJxd+Cx8Yd
LJKeVHBvYcrio+UfrRjNcVWS/Q+q07LXDLM3CPkkSwaxMbIXFU3F5mA4RizS789SUcLI69zQNGc4
h0RnUqzLE4mBvbRCazrrESH+2p3dviCESnGnj/Rz6VINLQ7PdAkmuoUbhFgE7j8qVB/99cw1aT0j
76ENpSwH6DkaAqgz+agQcC8j8yOzD2iT+FDyikYyqCsts0vDp0++3Zj4D33UDqBz6u7sOTntGEx0
XIljPq55VQYAgL9n8OXlwoydYkyjrYobQ2QMpcp7MrPxuGzqvrsySZohsk+cJdl/cBkjYlrXmAKe
zPtMwsusTAbEH4pARsuRf25rFfOgLuGbkVUK5frdCZK0IN9pfV7tWC8TW7QuTzr0+rHy/s+G3TLD
+ljiEgXd6R2IznmB/5DOUHAv2E2UVtQh+7Jx3yHY2GPghYECpims+X8Napk+mAQw1TochjQ6Gz5c
czBr3ARabYM9Kx7GmvAVbNrzWfMilALP6ODh0mdMyZVJijJAyMgDeJJzS63xmnbt12x5ZrH5upmq
I0+3nJhqlYqm/PfUcV5BhKZBC9YNprfXl8gFSu1sRoNPzPx6ApaUm7FGKADhlSgYtOv+ADiTeAHj
JEaX8HkhE1GAs6T5wm5OLCEhy16vesIW3IUG1mkJO9fQB7UC2Jhl6dCFAr7leiORiOzUCM2BDz3Z
sKOTNIEMR8kXMg019pMHU5cppWclvMUbM+W0ZMN8aIFWmrsDWTMk5jji6vqgl5Qaz7C8t1vGXpuv
aWq1mdlUOswCT2/JBstetZ5MiDdwTKkD8DmFqxJglTOVISl0eZDGhItgCTfabmY8i+qDHsZplxw9
gpvnSNUYa/dniPqcPE+j6gxiMgd9XdoEO0TOtY+tNWgwcnYrxQkW3fvFdMvg55KmINpr/5MH/pB6
dg6ncESjlV9kUTqPJae0EBwCTNB9b7kfNppKOg277iLgBJId0X6LJZNTfd4KwTFl98ct4NQejjYN
221oR86NaA4gZ8plz1MFr9SqbcZ5n/B2MP16h0uGyH0NUMsdkx/xxGDYJ8XSeyhkZ4Wki3EpyvGH
Rso6JOwUj0aRCgmAb8rG8GGYgiq8z5rxanI3dlqTEp9RaBUZrKqN0ZBL7irA6m9c5P/rmwMCRVXq
EaLTt2by7mSL/VLMAOF7cgEWdogAxTzcglDszBVATp1Kzy+N+SHIOloyn0Yn7kgp8uAcSdAMb19V
bznFV2t0ibBcgPOAHJepa1eHAVg1/YCVaypqrxtM9bShAzOROl/cA5t9XFBQYLIgIAxBhrNFi/od
gzQsnaa4Pz3zQiUNrBTHhnRNtp6tu7H1IBRvBcL0JxFRieNV3C7XDbznMUKi0gVoSDFbY1W8dFAx
/CTHnBFP6QT98mmFAF9p2DXKsCRlC4CKhh0cnUlmPj4SLr/7UtVRUJ1YyUKpFftfANTDwmw0U5U8
csJREAZv5P/XUTNnE1l2+SB1rkNXOb8xfnZ/I3p+mXewADMDz0vKWyh4S54R67L7CCViSGkM1zhJ
/OHn6XuzervAeO9g+jfZBfIrbi/eYaJafvlxLhQRgrJM6o0gviskivlzk5kzTUnIXhEfFFaD/tLf
b6d62tI+FAXJxOKEYjJgpBXplVIWcw4IpkqfyVHjvbzQZDwnPefaoX5AyZkOf3eaX76dyfCtFQ+R
qrMeXR7pWLoSwKrwIkHKROeIxk2a0g8QXj0QTuTSWLGwtkgBEL3gTEhED4CJgD2RKqm0DlKXofza
hloEvyEfJMKyErUmp9tCeHj+NTGHMhHCyrVSvYLFDdogknmpoJGxa7DONztjxFnKIkj45qlXk+w8
z862PiKKylneKDbPCtznU5l8ICJpuuiPFMcu/wmaYHkKOszfO8SeUoFUBngdmZDv6cLiaCzirxPc
uJSzdWGLZjjA10GqGSlpNPX2+k6JuoPe7TQ6TsLhbeLmw1mA7+YkqOXJXnHNDA63khhsCAzEISMU
tNN1UYljwAPIa466ihkb+jNZp9neS5lSHlTBRJTHsMT3EHzAf6T/1eKAoGdQz6Ndb+zYHsyaYWdL
u2mFfuUeNGwCe1vIN9fHgCV7sABqCG2KS/lz4j+m62OQ7JRoWfFRcdHsWLjseRqkPsSytuiY8ov/
M+FakDR9+FSmwoQXHd2EwLcl2maO6P2CORtmaeX7xChREOF9mUkGHvAjCk3irOimgFwT1X3sSvrS
Lo61Q4v5xplqIL+pGeaJS7QRHcpSdd+f8sW1CDwGEaa6p3oJ/6bJYBwWwieqLIZwFdi4Hsa3VQ/f
Afm33WUjUfdBRlaTPjkiI41cmEXVDdL2m++BCYnGl40pGKkq+rZt/bHNUNvMQz3atv7nlOwY/s4j
roWFHqTeUeV4aEGnTgK7sJisyXXPsG0aToHL0xPGpIpAJUAdb6KgVBm8urbB1pcux8tjr84MxG2q
siURuZ7gxsIjWFxBg6RAxi9rTuIYb02FWyLGXzFR8dgCPwhPU/SmaEE0gQh6o2sTQamhx2XKPCSF
M+9xKKD6h7ZcTPymsY7GYIgXWwBeKymfkI3/YQ7TJ2brZ7eClnhsBcGMjCuOde/O9OPXDi+CXMox
tZfmKLadpDbe1ZGvsyutjIMfsH9SaZfCvDnMEjvi01gtxzhZ2zR+ADrYQHWgIAai5UKkgNTCDO9J
yiOLcdloFy5JOgeLh0lJmTJVjtxBBPoiLmcQ0Eyff+E4EMWHVVEFD6PRsPk+S4BfattpGPQax4gC
s9X8WkSc1QOctzVKnULlkcLCE+E5Nwr1/Y8a4zir22wNxGa8aplbIugKkn68Tzany7x3vZ9rDiTU
6mZwAPKMPfJ1A3LhtmU9hpY08k1yDEZCwHartnbK+96rWxnBkXmExrd63wqBDLbU4UWoaQtVfI9Q
4lkeQntn7jTuqJAiyLcnesy3VN9oGVSKxxXNx1ZYw8XwEdXNN7dlCmER//XdZ6dj9V/2grBarMOq
xY1WpwYBlPXYKj6r9pJLwgH0deety0G01jQ0wPBkzh0jyO/j4qztuMWuNkGKyC2crQPh3tn1tV0G
qVqKguXkQ/NU86K6XJJ2KKlkgZnlgIELn5lNonnRKc22wWzIetBZrSB5/jDheaM1zj957gsMePFT
Zq30X1dCnQ0j3HvYfXyl9Ru/hsCeBPwWciCMzl6ihDn/sJGsK0iT22eThlzJDtK2XKknpkAL3XQB
zYzEpZ1FYpgj1WkXRlT0RgbCtBnKx/TerA2rvXoqEHIS97ffo8y3D7tAax5euro96s+wMBrHfkDW
+CPCwJ3U1i1htjO6hRTBxTey3ezSR2z+UN4/Bk6qJJEEFSdRWG2bAYXS4nK+ZQLCmdPbVYlA2Tmx
+yjGsoxuInvxUglqGNBsKTdF3e7Aq7JNdeQ1oBu6Dzoy1u7Df5kKigCH8esVxInWXqwTDGlrKT1i
PwDea0NUdSt6crsrK6c4FF6qeNGaxLFD6oK3yiogwaKxJnPV7sZqKz3VH0nRqpuAPQtG4qmMICGr
VJK25FfVyCwGmPlPLo3/7op2GuO+V5FyADYOmuADwmDEOm3DYlf6zNagl9q6Xo4cJOdSqpbxhcdi
lTwwtGa0LzJ3lIv1zGQNJSzZwiuKxIzSTG2t1HG167IewnyjeRRLP0epMsHbbqlBuQAG+r78Q3Yg
c7/uRJlkRDzEaMNEDZ6DNtR7fum3sniS8XKJ/DLnATt0TEazLq5fkgZBCwSnbIwTpOZFMxu96H0W
qOzR2+ac0XNX9s7OiikHN3xI8U4/YILkERuRtajf4pany8zzphvHc3PUNRWQw70xSuDRgcPKVKVX
1+50jLq84f+5rXLgtYgHAWRZf/KKu2x4vS6/WhDiY5Gg+9SX4w2sp//pPkD7X5Jx9zcZbl2M6BAb
Tm8TNotNDhJjdPCH/GnNkN0iRW77IgSPUcXuQZ3m2rR+ztxR3Dv+rNv11HNkP7fHe6dvNI4oc+3k
02hZYGmFizLTahjPDQGbmD+1MyRiTTbxifAKA5AwwF/LpMFHqtSbUqrKw3Bqyt+E6eraJeJQAybD
2FSNiyYbZw93RylUqg6/GPQcrJDOt8x6k6h/yH2HmJcOeuqMrxAx0f60U66flL4cXsIYb52C1z4H
YePoNkoyrrjZQb7WMH6ydNnoywJB7xI1HNPxfw5mfFZwwskcUg7zHE4Mjn/CyV2iEQzXlboo7jJl
RpV6LzdOjfbbij5JCPKUxIeihHDfCAZVoSE+/dc2AGVJCKw8scyajaLhdeb5ywu5Wl74FlRA8y3h
3Bz+dXZGDgjrBOw3czzMuBjkQnIxYFazgtb7hgatRXyOuNSo5Y73RQIV9gGGzzirKe2yke9Tskln
BMoKzmg5kRfJu+W+I3o88T1I8Nf/6VdJ2aFsKRiXu6RVZda9ipYcDzpCXPTP0O2TPrlUFOUew79t
paRSizO5xYa2y7Q4L1WSojfRqtjqE5MNPyZJbeSbGMQ+LHXG/BQX4zoCm8bvMq6OyPCED9RmTRfx
5nUu+3OAOKrfRgdXANJNFrxFQe439kBG2U50Rch5acEwBgLQLPYtNvKDMeoGC4GxdRabgQWOZVpC
9dCDM1LdinrdUt2aOxoycjBjkvokd/VmP/kBwo1qGh8XiQKTGy0IV2w+rXKNjY386yYbNySaudcq
x1WFOxp1oz6qoFc4niDChk0qS6V8hfqJCZs48Bj41qNOtdj3ktnlzQdAqsY/zoL0PKxKVlBTK+hx
n0DRcOm5NCrDDncjKfDpC8I6D5wQWhPZ0W9ei+iyluU89iAJKJuvFuLGkwp/ofCu6J5ebqquQGrE
21E6oulmNs0g2asar/b7BFdQ0h42myYlpzAlhWx0YoTtecvPgUgfBhbSS9Y6mKpwibMDSN8Ozssz
P/VxnZx8YF1PH4HdDY4oj1Tr0qYquMGtJkkyEN+bL4Oy8XHb+0+7BD1n0BJQpMWp4gOOjpH9+N7r
6H5cp9efFRcM5CGWUBAqD/rqTnDAapi4c89Xax43sZMDdrixbiDAK40PZ5p4nMhx9BbFEoYclg1J
yje4vR9K5xws247ysWJoDtd+P7ELPFtltWCPlkNJhukpv1qOB1uBTCDxgT/Z0kZfcIQS58rHTjcZ
ZSYwPI5fXJ2SSO6/RM1AbNNfmcfp3xDoN1vfYfdQ+2cNwVu/PUzxtNPJJkBiHS/IoPUYdb9C9HNn
ABUqQaAu6XSTW2gC414JsvFRypPpmrSsPkyvZjvGu47bP1LA2YR98211TPOpjlgLKu8a0h0ImgAw
IwOwFPNrbn06UpPMf935sdffqSJ0wozt5SmbcnPXSDdo6JAVcDU6xR7NqFUxiM+5o1DM2cBXxdBx
1QOt1gByOKkp6ZlYP9aVbrVdP6CT5l3sUyWY5xg63lAFX7krspUrojNs2UtZbKAkXhoPjh9VywEm
jn4yQU+ZTxqx/RZkdTbwWqk4Fleh8eTrd8ZL5XDMH3ARcPBq9xL2AfDxg+f5P6nE2w8Fuqp2Ykhz
TNCRzOzE/Jo3zmOl/9gdT8GJ+qn3Rf77qdnaGxAGmnkxi6Z5FTL8yLjoz/ssnzsGwnnF6VC8ktcV
iLRv3t3ovLQdH8uymcQJkWtfwNJ10gr1g5qq8yhJzqfabR3CNyzFyNSS0/qtIntrzO/vnYnqOHYv
1uMgcPuM3BvA1e1R0rKaYcQU12fqjUb59uj/sTLsWZdXGNRnsOqHo02wJE6160paZN4iYK5Zz8YU
2LJ+nXkzJzGRpkEr2grOG7FeMlzFiarmtvED2inX1SlXmHOBDKRp5u9kjwADP9Vw1x86Ihv2oCoc
7kLyyGC2pSSCMfgbAC6Xo9xwTZtyWu6vBnfGCaPNnrrv4ot2x5l5jKClUrg78j0tII6UyFOEYM1c
FIBdGamC7O0iPc8eY2IhXuPHLPPb4Uv5q0Z66dOnASqrGtMf/shfxGWBQqq9m/6wQIR0gZLjNhqt
0Pg7qXVg4rTk6pgEeO4CloL49weXPNR+/IJY2Qk1OZ+XWK33g54D3VUQVBATH4Qn4HF1Hk7Of1PJ
FQf3c3KubD+nyOJAiUjI1gEvJVfYBbQYuraegvw97tnESQkLQKm0Vi1e9IXl/v9YjeVIVrnUNNT8
1CIhsuYuFZW2HMYA/z3WfwIQKqbQRARntUvCLzjw3OPwwhOGv/IE+lywlbcHfP+GN8iK7SaWDSvh
m8+1DdHzA4ahSDRhjyC/jIsJc8EVYs0xrO4KmPHCj3rYN/jWtdogD93CoEq44/eaCuWreaU7EX31
fpMoo/WpxbjRQiwrZL0peaRdFpYZ3CC6ZrhoXJk3puDawVayypzxwmxpnCZO9qsesf9hfIY+2fN+
WO7INFYN6YUKKYe/YqZ4Yq9mcI8Uo6RirTwoyRqTpDWjyBQppmDERjtoJ1tIfuoBLyR1odduWyyb
XytGPJ1J2IHg5McBcalZWpuKQTWEqv2XYFDjANWpW+7uXGNMDlLqiCEZWBi43uTCtLzhMJYyEEPp
H6g7ehOXiGmkVd9MY1m8b1iPAZhO9i8LN7Ij3Xo9Hiu+WAXJ9mpdlG+2tk1+QkjFXzfXp5QqTpUt
EYj8dfHdjqDAizV2XB/XmNgHGVG4I2jxAGs0zWUnWJZpygC7efm5IHNnY6W3eamapsluliGM1Ev3
ACRB0BnDKyKQR1WhC2Iy2xNQANCd95oS8Fe0mkQwNfsAVuGBE9/N/4rnbAQxwkN4Vz9sQIsYUObV
rV8CmE1RCAi4no8j/kvNgvKOux5Pe2nhtUDaI5R2DuKqR3VKsWWTf/WwkLGlVJhirxYmoS/Dqa82
XIZa+Y03gp/upIFSoLDgbNBuPHEc9RF1TJSxtdU6mUT5PckVjWBSeFzQ/VoNu+cgeoAjLP9wxBNL
qFvNopnQoAK37d2Z9RYpEXMeOCoPbFVII0UcMBgXQnbwC2XuORdqN5a2WWbQTL1spcEDGkGEg97q
D7/JJBL9Jf4ptPNXaswmodPgs5BDjJk4L58XaOAZV5tvRcZ/Uzz7vaVVfHNB3KKVxjoGCWGBtiha
VMhat8ouwGjMF6UDaRD/59sQaObkkGZnAwDE1mnG8HYkWWfdWQt9SE8F9jfBFN55xISoq/Z8GqCo
JUJ/WXHjyTzE5txpqjru39PKz/tOTMeagfACK74qHvsUiLewYRYatkJuSfXQTBD/lvS5o40ZpXuE
ptCXbMno1tPaVniSv67tdOA4ImfKlPw/27LTfycpHXdmsI0SgFz4kiWX1jRckAzIHh+FYliZhNpn
SIsD/DJAKmN30i7TI1azOgodh9t8Iud6lB0JQxHaln2khDiG04xMg8O4pmY3dEfjJDsym+2i/AHZ
uBpjsKzXu6ZQJ2Fiqi2L0S+aptXbeN0Lh99thwtIIok/QuMYYIejX1EEKYpRUz/f3+2VvrGG/Tbg
zOpB05kBzo8rd5L7by9+fJ9/u7X4OF4s4XXbGYzpH0C/JRrFJTBmOXRG6miISNUCoViGAEoIf/o2
IdNZjBEGz16XGdwz/YCimTlDO3r4yN5t4OuWdrCbIXKuvTeEUAcuOeWuBGveOVRNTpRdRvzxqfNz
nR7ZBpTo7mlKxweEaC3HqlB7F6MJ9dk795Hc438Av+v7VB2Oz5Q+Bz0vf0QCNU4p4TVcvcjQtTJz
OSlFbXOPn6QAwNB5ldoN98eWKn7UtmcENm5BLTEUvCOYwhQT/B45ajvokDnwg4JnDA5xLQEfGXdD
FZaxelB7QCsmxJ3iJWGcnXgTlS5YPqJwSiHzjfNB9VsRs946ZUnekYArIfm+0cNZseUIAyJvngVB
/LTDbcLLF4xGDhK+6Bjpq8rS0P5Bu+Y7JjBLp/I/TGWhxvznFpO5OgLnmyWt/4IEFOL+Us74sinu
N/7ls3hs6sUH1MIm2QLnIUvdeWl0fxK+scJcTsWecbnVq54M9NmPCAVEWt0pwzTH1GKqsy7I7Fic
dlLTC1EY4MgN2y3OTjGkQwXFNW6qSUAnXP9V20v4FVhpPoatrCS0J6DDVLqotU3MQyvzZPil+OyS
Qpx9YwheKhDm3Rhcx/orTiWx3wrTD/8qpp53zjCUGN2bQ6sDkGlafh5vuUAqkZNjnZPRcw0QmSSj
1MQQ44ufxP81tA3BXxYi/tRfxEXREGZQKrm73gSAKbaQ7Cjaalp+v8+X5eTj9836jjUMlHEQuXj6
jy20yj+OF0iSgNVp8xuzkQMwuibt86qI4GSYUVyjL0v6vZdQyDTRCBsP0q3ESB2WZvmfyw1hSN9Q
zmuUkIAWEnK+c5Y864+NPcJSSLULX9n6ON7wTeu0uV5sHZ0nojBgj1utiGf6oawHiE0OLYtdT2UJ
xAIiduwxR2FnhJaXgyKPuPrmzoDeiLJXXBtaNyq+IhaFmT0SO5ZQ9FIYNi1MSzNz/uCGxJ1amRjY
ItNzne2tdFj6HpKAJyLxT8hWv8LTk1G7WiaKrrP/S9jbUtxFN0CV1l+IpB0mjc6ndcnwEW5dalOk
d1W2x3/S8F79W1q10tPR7EdFBAxf8R51fUAePJVwBleMGXGyKLJpe/689QdS9/F2JxNP/QvjHgaQ
67OWSt4+nCPaylLBrbLwVHNkDM4ELOD/NvE/ZqHB1jIcEWfyOa/1BEqS9okBxjESGYsT5CGSG3TN
xhMoS/86OjoneU1KvCiv+W9GfEBjR8umb+jzY1YMOetRgaav1knTW5rLIngOti3WuyFQg/u7XUSz
K4ozE0jHflA4wadNAKXrqIdn8nGM3ZuOw/kzKBnBsw3fUdqBJUXwpnWUPGX1UhejuvNPExwNctE5
V5DohbVkLMGMLX4+kBA/H+X4PGRj5dC3sJMovjj+5jGQjTfjbm95Alh8dWvGU5cvFRcBkznuUnp3
Gp7a/QsB/RF8A7JxKCr5FaGY2j04QmBHXogeDOBpRvzNLw8clt8wqIrVoqIUkJtTycxpZz7A5Urq
9K5xd6vJG6nHojDsuySQRJqTl/+o3X64XnyB4ZgsmwnkmMdETlj1X7nIfCObHnP2t/MS2M6Zyjgo
kBpApPmV4brZKgxl7xaKYGoOvHqItF82gLC1eJZYDo83BFpEcA5hoWUzbzYc3a++KE4Fikb2n9lS
MgN/Bku2f75pE4xqi1CfvHUzEe/OwIHbv4rrNdOwExhWivEXUxKqDp8nAXfMMgHDi3khDvNHrk7u
MCQl98U4tk8yAOgZI+q0YltgObnvTgWUTeGfYrG1RmKWGa3hKVmAQ/R0al2MzrSMTpdvppQF2/bZ
nbHryLsYUNnPNKR1ztwruuwjtzirzUvq3nAkjycRVBagldghHoWeUNGuVxjzdvGegFBc7URktEu3
WdWttFcICZiSSjiaqOgL/BfAuDUmDfsbD2tpbnyT7e+HYbIgizi7oMkQmnHvFYMU7/bALOPy8HDZ
HkyXgTNc7In9Kzd9848FfRf+9p03VPuOTip2s0YbM9eL8b2z4qitH3QsghD5EiLNE23qSYIuj0rU
iCU0xinQoInXoXqod57qPkRQvyFNfq4+RzqrbVIRw5LUdkPVKoFQE21WjmxVpVZQ9MZ5XK+WYNFq
LjAJs0OV1E4loIoZf0Qho0lgGJnIlMZFufdThmdomwfxajQqrdQ2RC2ej7FwSYVcvJMZvqfzCUtz
/uXg4o9/ukfXlFvNDfYNIKyHitJeDyySrJnIulkQGw79sSAh8kFiYnfsjO5eZqlP2by5tdt9JxfB
ZV1b2WXy7adCySxdEyYru6EC+AdxPk4qtYVuvvfQLz76ZiacQ8wn/EoUhhu1Bc6iS3Z9IoXEQ9j4
twxoT9Z/UtikDIbJgmJsctUZ1XfxQX7pggUw5YR+VaOhgbWIxGTh+S2KkVemQRA512MLVxaeICsm
OZ6ThfaWTO+XZ2SJjmLxyB/77Ra2ES7cZLoMLvIonO/wZki52i03hZw8xBTuGsMkpYdj4O9Ja/ok
SyuehCgAXE14dnqKWUefX7O8W88WND+EJYqJ3EyztiZrYu9aQNzM9j4Wvilc+DHQPpZ2P4Bv49TQ
JnCX8BtV+NtR+s019TAy6usKjE3EUmaeJlGZd2yblrDnJ0kGIjtb37bXXmy3LC5LAsWRtvObciVz
yyKLbqgOfuR4r/czctS6C5r/e1KNqPuo7Mf99X+6TLXUTZDyWtUC3GPapljG/3bkK+hmkRBQrT1I
8QUeShUUDvc/CZBAQrc49fU4VtaNuMqKAVRUY4fDHKeOAILR9V8AY0jE9zqSPQh8tmkHm0oi8u49
aEyFMUQrlvEsFuE1pvNzJit4wk+nM1XlTqlg2ttZEd9+jfh5evDBBlODhW1/P518Yoou1G3OlF2y
JlZupaakNPLrAhcKZVy3/HgKfucbSA24yKwI1qI9EOW0ZblOOdF6qsOeStKEkITO5pb+Q2i1pMWx
Km5CgkJblEvtzWSF5FKGlOqjxDoLRa5fglcLjGNRLg06luIeZBCmvXLr4iG3w5cnR3jNHyWT36+z
zsPdNcAspq4JJnaPZhMQQlI/jwLyC/4SXdxOzgM5t6Lh6vlaBZeORoFSZD28i8uIucFQaQDw8c8g
4bcF/a0bdFEvQQF3p0uFZ9Qu/0O5039niLFTcabXnzX+sp8Eh1luCE6Ilsgv6VAhDZXROqQ+8TvJ
fpX/9lGZw4wtxqOX6P2SMgor3ZEzUhHNUXlkiT7rmRzuZs3HpiL7ZRQqZmAf/Bui8D0l5njYPLHy
Dp63EcfvdSyh2Y2eXSLrBS1Mcoj3nE0VLIyrtyxZ+xTw9m0MlAivsh1gR9CtvLxt5gvcK+M5hFAU
7Gw7dXWGBU10jzjGfAlV9p/+qXsh+Kd5gvRare+0YyeuUMrZ2sUnr9Fua93JW+O8+6LhCJxS3OfX
KP1dD6cpatRQMHcy5QWQI0FLWvvfmdKxN3pBR6SjWAut3g4SQpEFSTeKss5cVVIrDA3U8geFPSGK
3KJ4KCQxB0ZiNVA8pg1g773ibf2EF2FOi8jL1LPkdXRj85O4rIA3TRkdPYm1H9xU9QLG5Myx+gkp
6ph33wFNla4qsqAZHBrAfK0RwEtbcSZ92/bfl0wuumLAufHbaqbyGd8XG8VtxrU229ZtZqNN7Ody
i8nS4mIYU8RqKTyTG/vthe4svERtJDT4fJN28okIhLySv6eE/1480IyGyptPxeTEiW1uzAC+Il3k
FE3B/0bmGHOJf4AuPl9Gdlxq6rgrtE0FSy5CX6fPQNHVCRlPAD1NzJCpuG6Nvi0Ra5xVz5izmrOX
OOnuP0R8GDH6/sLeJRn1FUU9A8mxCniXpabaLSUaoxa7kqjMxXeI2JcTXT+XL2zOs1BCBTi++dRh
0iRMEfFW7QP7v5Z1sqTyiNAi7p/k8AVPhoQcMnH8hn0mMXadYNhZEE4FXgYpPSu01lia1tx3L7aJ
ydXAie4jAs94ty6vIlJsZnof6SAAHh6vrx1tLAKBOWmlKI0dIqqY79scsK3qARPX1x3OlPG3uLdg
PyomX+DXmxtGBJQKDb5lUetQAczngME0ZyAzjHPEN52mIzF+ldIbsGX58LVyTB+s3z28uApKc93S
XL9x/VdMix1qYaooG+a0z25MO5FXbhk2OUv0OPeCyqjEJHleX452UM037DgdZE9UNmaqMoy27alt
ZJ3nkAWXupYrXk+BDRfMws1pgBfeKCazuyzXbnjb+cgbawWo6Wvr5CJy7t7E8uznTR+h5cup/V77
VrVm3gGH3iDZU4cQaBw8q+Dt2INgUaWbZoO8+JzXuBNwGcvtC2IX9eVGzrBGd/RtxmRh+HNaJ9kS
5sJ/xgO8FeoESj6R/pBbQkMJO3/9TUmLopZLh33AVGeaALuaMD41mXlc6pifmnjmCwr1clrCLAwG
iDSmOGU4LaPXzw0FPDHop7BNbc8lnSRlGxDuKdBCqC2HoRl4WGc2tGe9ySAkAdhL65zivQmsTDAv
rxTt6x+NoIL9GBi7u4qEQ5bsJ1zrWq4lpqWmoH3hP5m5Vh8609LGD2/ZjNYcjMBiWR2hlkYG/ShC
XZ1n1FV/IQ592xGHqAh8d7qSCBgj+JwIS+cC9ZncP/96x8uZt5v4VZB2sgBTpu/T9bNhjcFVW7A6
7n6oh9ozlrnX6JWpJgOQjdxVzKkReN1ewLqFvKRpH07+oQYc4ovFGVOXfUE5KZ+mQt3B4r/2lIY2
loo7ApCmrdeFzfz01BiGniGm5fkoZK4H7cc65M6Ag/nNzV7nP+eMhk5aOXrD2MVn/BpisuUnYiPc
P2U/pLoaHQ5HqKx+qzktdiznJwHVygnNw76pAHDHMDEbSvoH3qEFxdE0bPm9WQqWGnAgzXb5XHQg
N4Ddg7HpV4LEmQgDU9avhHRv1BjUDvSoVnH3CV9B923r/aiw54htXL/fD9FeSKd403dw+iHCAc7C
ntfXaMxj7vhMAL3wIiApggyZM6HdGGyy6m/4q94HhGxjSX71bvftD9rfbkVmQcxJeUX0NnsYuTWy
AvilqXaCsOQniAMNbCOGGY8FGE6c55WV2HdEely37WL8EdqMXo/x1lraGI62H3FR4SPx0ja0RVly
6xq0fqQFdWkpiJRY6YXjVJNbOwqSIHxAsu7UXr8N7Mww4LvQImHHjU2UixoAfA8ecUo3jLh0fsz1
1+Rjg/drbMhfdfSGNAsKIXHobWw+CX2j2IQyFOyOtn2jPAPCCFlu5nUVdngOr6vYh8XLmGnv2EHu
E/txuhv1skMPkCrEsZbrl8Aszpe2ZqUDF1zITcISlS4tLOABYfbEnu0BeloeekvhiIXiPkS340FQ
ty6pLjkL60QvOIhYyEzJozHyZBxd1XCPJjzMfE1w3ocKuIqeGeWkpvYi+KgsKszDYguINB5zCDuC
KnLunXRM0GmIlFWdq6Z3hjoxdcqVSqfZ4Le2JDxYPTbjnM2p9w5QN3L8t9Rz3S5xxIWL+ix4p5A0
t3cUxJVgPOU/1k52ajfpIV4Zgimn8SZ/ISm6jzH83vbfcWRq5YvFlEm7X2G9MErLEiWHTwa9aw4L
AML1GINKzzwlbD0Qc6AEtPaAminLhj/zVd9U2X0lBwzHKA8ekj+jgTQcCheOtlCuvNB4FmJd7qbe
bcnkcAup67PJnvTnAyekEinOulL5iNNPJzrgaHl/Mj1rcGrk9Y/FcOQQ8m53zNwB5zHVZW0DwGtU
ub49mYi0aG2t43i9WP8A0maHT9fMxtovRdyUnrzP3GmRvf8FfX4TvDR203ckij2B+3m7I4Lnc7aj
XcL8OVgXNtu87ERrl60m8S1rdWe1MC/NvqWgLpdiAi95qTDSOMurp1+5dvVsCskvhymPdFYOP/yQ
nDcKH9ljH76epjlB9Ie84RC6SYKdg3ssk2b2yTaIYm2XwSVMyOOPQN0cY/qrO9CwyGHzyQnzMY5k
8CH113oo6exnU/XIeOBouaP4/MQ+SiSQrQxvserFH5nQyHu4rZtafHt2BZPgaAdljeLECAEAoYGv
CXEpeFXyaGL18RSf3noki5Oab7ufCWCrMCIwfCg9zkE3+PHrnHJ1HdhniIOs5R+Zt2mzSxAif25S
/oTF47YgRNpCzuH86MN4CtmrTd5eoya+2CerZGZokT5NtshxQ399oLDAeVu/y67zolO+Mei4b4Ki
KhC3vbZ+lq4HyeFEY1eZj1YyjRuRtcSVxn0B+1mgkuYqxrfjA9wE0aMJ6JlZiThATZSsh5moQrVh
F6ZHPk/zCyI9EYQJye3EqMedr2kZnxJmclxEq5EfswlEiPzaXepUt2jycRB6tSczyPeXU8YLdMrW
0wflnYSsBamyJzgp0A6m5fxmDvhfFkvFEUWyV5pdLb0atGWevUmiXoeqtQlKOitdRen8jK0Q8WHB
DGFExppSffeh2hUeWnWIa66sGmp4Rx5mnVdpRJihyq17qqoR3RisHijAYGxy2uB8Fr2QtbX5F5rd
4IB3/NmaR+N0mrEmrML+nyI+cy9F8CD58TPhqvfcT5VV4fgvx7F6fXd02SEy1m+pwSfpWGi4f5u3
mpMqE3hcLQQJys966Xjd3gg770L2kqZPnF/9U+Opqwum1Fc7jIElib+gXwZQIdL42Ud6VjL+bVx9
aNi4Gfni1BWCZk9BWdhOr0H9flGp/YP1MaGFwoY5zN1bE2In3HXl9AyuTz161+j8ksJRCujeZT5Q
s36ef8tKp0G3MFRzg1ZkjNC51WqQRtrBSAdTBHIxbqIJp82UqZ3GMAmcoNYCSV3K0oOACQjNx/Ap
Un2/mOt4H43xkab3LxRIjUpzbj1x8bZw2urYCsQgUt34I9qSRxtWNx/qy9XgWExXlXKSPrzx5M7+
Ccdrez77kJF6AJHFpIqqBhdCmS5T6nzcbv9l8nzp2zezp1gs/qDM1kBtxyTRJi9WtbMZzcJvle/J
KqX19K07Q0Wf3mK3vk2ZJ/aqT6UlxxlLC7tyiyKfrn9XRrpbAHZmBMqEmP/CGxLqB1xYliHFCrzy
Rb7jkoB8POlClAQvrAhcB0Tk5A5IuOMvAgG7u9E245pkUknOTJttB/lwXL1jSd+gjPoR6faO3EOH
JJkvI3YDPNTyElF+iETylYCZ0rc1dRaOi9RXO1xyc+3YP4mTgR+NYzg7Os1pM3b8Ifl0h9iF/Hn0
cNRmwV6hXkWcRYIDQ3voGgqVyUM+aWJOcsMGkFbqv9APP152fmZpvKidUI9xDp99vPV/Lu05123T
omGG0Z41ABll79aEHIHuH8qC1yjv6WO2EnDzejI2aqcIs4y7KV8eUf9v13QMkdh4s6/zSL7xBbKH
a6hoxg3Nos8sB4JER/KNk1tTgLn8gc/O1H1YjEzu2c9ZtoVxwmQYeWGTsI57It3tethu+51pDzHS
94FO0hvXTBz0+BEZK7HhN3MiGB3L/GVgY7pEQjzkZKdm75kTVk4PXBoq7BO4pW+BeEvdbnMx97lm
fYulYnN3yj/IXrjedaRjE9FtCARV+OC3HkZO50DYqq41cpnX/lmbTXkggIxpWBI3xOeulzHX/N1c
AwH0tB6waRq8iO7xoZJYZLp5jU1mTQexV2gP0rrrJyihrkxvn38jh42us0oHFA6vLWot1HPIoplT
Ns2nqgygEBmxeUs4Hx5T1efueUAoVfB0/wOkvPtGvNPd+6YBAviGQBgFc5KenGD0vR3EoJfJzLjt
+fi6EFXOVrGbFGzsDXBTu8/kfdm/0k9bp6FeUBa9ZpnmKum8Dl6ES/kjc9eh0KgjZC18xwOy7NCF
BDc64Y8KrL1ss2Dn8EKgKwFsCEZ4fkod2gLL5Vtk/yElRs9CxQToeidHtQQGSX6cK5cbqevPkT4s
NnYgSUCQs3WG/+OUg1W5VKovvR/jIoZQjLvOj/ncy+SVVqXU8fZPquJXVyW9iY9/dLmjnB3GCDCg
m/jQ7XCSgYaFDSsf1KR7PVQAB4xDx2W7GH3G+F0MYKwQPotTIpsfJwUfLj6IkOwQ0YowAu3g2hwG
9RT/9cm3JWN5FaNOh3uOGZLEa87YrbdIT+PxM24n1QUEplbwy5Bzc7RNYAvf7AzwGbfrWzQtK6s7
Zrrd130JA0bqVjN71/xc1gLQx3twDixjF1LVZRrWbKuKQ1soE9Sqrn8RP+q5APenn9J5GJfF5M1u
iGwsOeDkd1FUeaJqN4WD6AmibCNCKyoPQ9cx7GXToKE75NL10iemla0kys8MX+ZWJM0kxVQCFfv+
0V3O+U/vwIJu+SWm3CLBX3EElI4GssAzf8Cy/HwXrKxh2IWkj/xr6TdjgRkar2nHlOHRtQxJAKy9
VfIaolITHuzbZX5HnboPoR97qGNRw3C0EHn7viy/zRhLz/bABTDWRlrzIvvPbjPrlla+OkdkP4W3
LnL/N3hjDHWR/O+LaqeTILFOotA61Ps8gjEa3dVxa6PNs6BcPa9eviUQALumWu836C/XQiIo4utj
Xl0kxefsXPBqNH/Gc5UIKqvRadgtiBS0vG11jO5bVGCTBIcjl3H5bBL6a5FmUN8DIqhw+5C8S/2A
4c8B3HDWqEGAF7qWU1Vpyq4Gc8Xw/yUtMkC/ExZFW2Uhn5FvrKF8mlAAYY4Xls2zfCNdKp7PDvBq
ESeqF++GwnGDUs80MvIgr2CcvaxvOeNHcotya9w+dJa1EOpz8k1xrBz8phknGBuv0gpHWjkOQMWe
nCju9kxg+wEDm6tpoEYqcz26BgfEHPEx6KtAQTMNpTlV1ruIBFjHNrb4xuDMT8Tzj68vX3TsDPVB
jE3JTRFpq4yElmYVPlQl9k/OuTl9RMgAXUQ0oQgGb/jPvrLO7ao6wCbN0vVS/jXLhAry70Whsipg
ig4l78G2q+YYZ1i+h4joNP+n0LjhH4e4FYZE96MD8cAOIkGoIAypYSweC9dhf+qbyaTPtvBzvseX
FPB6j+sDj/6oTTSQ1HEYvnW/VO84rcorPAWdlCKjfRsSTu9wxa6Wuc8oTuhozD2o2vku+Xjgp6Gs
FpLd5QQTSZ7ASrpReR74N5fcK+4PVBfY9TYEi29q3qDo5Ib4q+riWuTgEvqVftEy1//ZZ77uSKfI
eH1NrfQbSgYC7nXS3kT9a6Ly746HKRrsGzxNL6rGBK3NncyX7uptVb+fNA+JbYHJMSutAbhbCKHD
K/htI+OfKp/rD7k+CIKu1s8NiUAQ3bPm2S7fIl2/cKmQM1ydJakxrrPi5yGhK0zQutcjlsfOZs7K
oSD79wmXodtnQb9XIeDGLvMYCAE+F8kfkpLc+bNLKrEy2yaA6Wbjbgga3Pn8u/SYoDTXUokYqodu
OPq9vEhHa17zJlyH86zBhEULgqb8BvNP/02hBYlLEgCDMJ+bNnj9bUBBeYCgdyyJ/XDIox7VBbb+
yf5yHXDYyQqdNIXpSvG+hff9JGhTidYi9DmSC9OlPQCyyZTOUFZGrsi3ub76kJqYbOk50Hv6daNm
mwCfAOKFL9jLjBKMvrlj//teMjytJtveJcBuibNWWW/koCleSdThDzWEQeXYg5YNRf75H+KTj7TW
5SblzwUg5qIfnyiqu8EqB5GGjdZIPdi6z4XD18qaBLDLvJy0zbLmOON4ztCox0KF2LS18iSgMMJD
hqGTyNRFVjZ8eVvVSIdZRwu6UGJ46BclJPEoYapr9YXYLx8OZnz27qgcuAOjrCd5tF3sCqcQyVRq
2Ohit3C+0FCUZxzxlhjG/EEwQ+7gysdRFaTA9XhQr5uOO/WwBWk4i8sxNdmMqZXtw4NGyuQrAs30
p3lIaiz0D9Njj9LcYKZ7I4BHkevINPWd731G2YycxeunKI6l2BpjSbvSq/z8o/b9bzSWc8uANh1p
KrRrvggi/x5a3rhYmCuMo/K037/2BM4OyrXR9VPRsSSGovieAFp7NBCHqJoiPXg/TIWOHB3e/Pg3
Yx6yGVBXRLrR5ZeAbNsX5GS8vVLRKU3TSKVa2KvGILw40z6wVtayhYw8JGNF7SndN2V9Dd/tVDOr
nb93axOoq2hfx8xpunFZ12LiOEKoDT7LCy268iRhFXbYra4CyYIzLS7IDuv41Sf1iHNWtkYAR6QS
DID5BppzXn0/JkzNLVLNk5hlnzqvu7iyriXtUTKTAWvyOet+TObSpDOC4cKwsGKpeUIvYI1WID8Y
05PVn4BCOQoR0AZ6k9Im6AHkp2VdIBw8RplQl48CEthcTWnydrYtXkevRnaI8tkq8HW5RPUi2cAE
Muq/kBMBHOcg2JQuuiS4atEvHqTCagQhOrPBI8SWf4mFRuy5X8IwsEuI+3BgU0re1m7jLwPxYtKn
OnNRQ9e+vDQYxvoJdvITMRwZK17gxOoz8yMndR2UjcEAVSrUvwoSwK7M9d4GFTuvSmYZcrvkotqu
vPygU5H7CZG6XN/vFCTx4MET9XLlj807iMKi2us3zk6yTDWpDY+szg2mCqEXe6u6xE/rDCbKU5oY
RdJt6KSD6CtOq+ifD8UZVFgFJ3f6FhOX5Hygz1c4jI82w21ay+lfhayHLgsRnyqAcvnhH8KrFsNH
cMlmk/1yXdRATW4Wg9Nsd3kr4YDkWrJ+ErInWlEz7Y4SdU1RvC+D0ciiGW62xvU9xKPdDfvi1hfY
OA8UdgpifvbEZnfNjSaBHRiNz5GumYjmDYkOrYoQp7/mARsyVpxR4PcwJycp9RBtilfBGBhQeZVZ
crZJUThOHXt9Bb5oqXhBbjm81F4LM8OaeFPMbBypmOaqwjR/C7ThEAPEVOIjMfWg91SrxN2dU5sF
pLWRYy0b9QQTwdV4CENnySuXM46ekihVAGDweYnosWGNqK6YQ0XuVr+0TXcTbPdSWOQtmLltTgIM
d0N7QlsVWLToQj0oBlPJ35VE9JcJfPRqr1r5XmbyL7shC9HXowu0sAa/a6OvP4N44Qb5s/+5ZV+9
2Z1hRhPP4TiBjU8rd7zpMlWOCjAaHN6rjruSrAStQAp9V9snY+yYmE2sHljvFi6Fa1jxaJSDgMnF
6uIH509IkO/hFadZkmxnWKrZiKEWB6gKFzW20wlbZalbsnJJwtl6zcTYBp0JRTTwQgxuBMcHaAln
Pvq1PXKdK3n0c3pfO5t9dbI4TQAMpjScmsv4b/n6ukpZfApymQrqMFRz6z4Hn+muge69yzWMKDud
M7wqXslYobtNnt3kfhMSDs/CbtiZp0Uhq+YH/2dUaLNSnJov1VxDRzbOcB2M9YiKvTzmEhSIuOHO
TPb7p2i7oSpwNiO5Z7U12uFT3hOFIcbEXe5iD17ys+mgPiKjGI+TwUtTHkgtm7wCscWrFgr8EuBa
NGzlUnZaYCSxECIjJlCtgcUDucg7+VmThoTRmRnRqaFNcadlmwEWSadz8R897a9ylD9jD82S+Sdu
tiP4e9mRkcvdy+ukng+df1FVoUgNyKzYn0OwqtwKjzXOkDfZGXuFhDfyXK9ujwh/H1V8ts7qoSnu
on0gLW7xifnDbqy7CHgVgmRZBVfKXzb1zvlVYS0SQc8/Us5jS0bjkKF2XrNTxe5DJ/mW1dxiWUda
FZ8UinMCVhNpBDefFBgI7+7125wO2VTgt0/K4U//z+clWV0TUCCxtDQtAHqAT0PL9q9d+X+PJIU2
zNcBLY5+vGfAx82++WYdQYBHZsGXN7h8VTiP/ZToYoNk1vi3Kak8eIOEbAB7p3FB8W8JWfkI8dAp
n2UfVjXFkRVPqLfY1Gsl/8pSQX1qoKm8wLfkkPo/osM/g0m7ZrNN67/bNynqk4eAUjQ1q0vrVKpr
tDqpj+HAT5xEncdtHflxLORAaeQ72WWwcbwierzKRKbMbVBnU4W6A3eF8DTs7Fl1rmRjKbbcKknZ
iRXHpMPtcTIaX6C4hezki+7WrUg4bUCgsjRkpGaO9WmqIl75Q2lk5LsRY/8h01umHH1ui8SqGq4d
2zOCAtasN7TuEgZuyGQBEDE1Me5LoYe0LHrXMjcI3nQWLAejxNXRethRhhsehauVqUOhg2MVnNgX
/IEMYu66RfWhm11OP5WCJf2OgmcGoZzmNFNjjATfrou1AO8GlKCBuyWhqN+qPl06PvtpL5PjfdjA
m3DDaxeQ2XNtOq/fVfJUQ8VQSKug1b/vTS7w7+WABc1ohD+bn/1RJBGd8QY73qKx1sJNHuZDCwpU
HLRVo3XdcicM5jhbuxyM7UxuUvIBEfhxtETWri1I2LGNAIGeuT6rQ3FJWMi2bIaxhrQqrBUW5tNs
Lubth3mZwHRoX7dDrSJ7VQwzw2qXUvM5MK+0E11JKXmkWz+TSQd5X+e7YjzF3UdzBIlM7zx36iEJ
tvI/wUH0emCY3uZjOCAMEzN6KeWplORwfBYJx4+bTVwD5P2/DZiWEpO/h4C7FEsEtRpx0OGZttRE
P/fuIq4ZxxwfSWo+zDWyUn7r5hlV09BUvpyKMd+noDqx2gMWTTUV4bpLpLBomlybJCxVuvkOj3v+
UBxxPX1p8yIL/rBQ2wFSOdrMHHKWR4qZOOCbQEqJVnRBTLqAPiJVXXg4LReSKz9KPmY2ku5wItbF
lleUZhx6yY7NkUlBBYNc9i7d/F57cWphwaFGuxslIDixXyxSACXUlVpatS/bPKv5Pusz1hGaUznn
enc/TePMYSyQ7YqPKpU3QkWVbXI9N7SjqpTWd6Z34zIhcCOidLn2mvHJ6mFCko2HZhKf/8Yq4DWw
hc+ftO7xKnrmRjElHv5GCuWhShArXOFD4rmDhAmCVmY2/i506hfBSO1rMITB7aib6iNCsvoZihtV
nYCnNT4fee1xpxe+WxKVC3ZK7kBHCnDwtfhcFLBD0K7Q+Sgm/PdFACnrSx2lHXJ0mVB8wNJnkZtf
BnqPxICkh/0IiJaeg/iQPe+ua4BmiWldKBkPzhAyAb1h5OwcY8a2h6dOz5LMD3bRzrY5gSS1I3Om
I6PnrWNV49iY0h+TGAHuK6b8eYL29m9sN7IHPWmJH1E4m+lUofN2fkj+8eMr0dqfBtENsDbhIWi+
e9Vqzj+VbKiFhRx0urAOrqZod9XUcC1TwqV67ZEMmlK6k65OUNcprvwfIWxK6lwuIaab8jItH8Hf
x2J0Tr8U4XpckROo/Jaw4ydQax9oEaCL/5NZ0luqE2p2NsosXm3ylkyMgeY8yMZK314Zg/x3edKP
w3pIbES03jadNaHvQHrnVvK/vH8OE2p0SrOLxDA26sIqDZl0L84ZAyS/3aNjCEExCsJrQcbjn0S/
KbUa0S6H+YUb/525U3R6Az12UWBakk1Gh7h8uWgjC633oco1EP2x+jhJhtw2n4SueAhjWWPuORnj
GE522zCnUhZuV+mfMKgXr8fKZ92FOwNTBIca9igSSG3D239JR1XKhaz82PvVpWd6tUhGhVjKmo9S
f/uuK/zrzT8wvwUoLUVu2rlOkCWupl76MLid/aIga+Vque7W0AVWXT6UDGFA7Erx4JT7IyY3+jBl
Sc6Sa9WwasIkhgRCMi6zO9mXTveODrAvvHcq0P4oD0xMjkEFEorDhhxDXEfBt6o9FFstrYemGDa+
A18F1UdVMwVcPgrvSo1dmSl8J6xr5tp4jVtXS5LQaQXDMagcvr/8k6ZVBCtgufV9RDlxqJjJImsA
iKZ/EZb+bQktv1rAk2n8lqfzHUCps9euMEimG0hBsBxtVQv0TViBFP4PGpTtYZzFlaVVrHuiH0vT
BV3wLi0gJ7MNC7KoxOcfu4PWz/nMcJjPxhZyOnbq5Z8ad2hE4VpR6PYt53UQExvntvM9iGFk19p9
rqDZ6CciQYevXn2mqR75ZNUbMJXNg9zo/tw8tB3nW5wotNhf1r1HxP2Ae2AXmTKS/NClvYtnAaW9
bvfUtMtVKuTjdntif+dP0aqRDEVZQRlwQY9WSgUhSc8SArJawGri6JjCB0ZoehRvEEs+g1B1IdWZ
eBjRKyx8h9mSuhLInoe+VN8eJf8LeaLpQmtxs+eemXiRjtySvF9Et9Qn9Uo3mqTVVqYR9csdZE9z
4TKiVyDLNWxYVm3RTJrgZMo/AKUa/53oI9l5gpYUcHUJ53XnsjyIn/ucxV/EDzcJrkOo3NVsr1Fe
P1mpbTyMfhzSSKHxvTAOglRAlqcyeIf+6zLfx5HHDCUOUqscBECV+4uV/QKfCk6n50Y0RcJzjBGq
pgLKR0s4owzcl2pX+UDF6HtKcRK2jRGAvDCqahHKy4MSWpM7f2fKqt4Bn4lu09r1VO53KaJdbSJ1
4iWUK7Npy15celwHIyXtB5uUsY5+bCl35g7cOTFgdWl/ayfI9KsUolaeN6lcNAjR9jXu+bFjyQ0+
6+YXxjFV2bI/IK4x3j0Bzwh0qy3Xvo2jtWMucV/tHu/s8rUcCEobdsbX48DgT7o0XBBez9CKrMQk
yKrDE445qgd2LB91M7XlxUByXl+3TlnD85x10nd+ftMPBcfyVj1UEQIe0z6X7+owdMyi6ckGkprD
6HGhkvjMuiuKj0ogcJNQSy51QN13+7MKl2079kno+zlQ+kg6YAjpLVvMbF4RJv2iwbpKIVMtLev4
Wu8AnsqTMuGLeAOcuMa9EDK5tjP56VrojNq89qcDsXnOqLdgG4Yn9hFEzJ9ze08r3/h/r7I0Fik/
SLwdjlhgpzQesrKVFw8gE0ZIlEQLhYmLjiKVpt2raKLHoUYAYzkAtxLIrM/9kjXusdQQ34iP77Dk
G4wU3tFUiFgX4iSgASlRoa9PmHvAFdPRSAqYc7kOBjqcbUcFHiO/dA0lSbabWoXm6T48KTmn4m+2
OaK9cHJqjCs0Dipg/id2UCRedGzvqDC9TfWKoQ/Qn3cXoj3NFBnqO/NfrtpmHm6O2ra1AvYR5GDP
OR6as1oInPYpPbo+YJJo9UPnfhFLKN9WFk01hE0yETTNysbwxwBosPLnvRWFmKntvuc+NfGjqe37
EF2l0M/WaV9gIcTBN771l/7M1bTxWds+d/MFxdIV18EFMw7blFy72zHwsiOpycpD759ctR8/X1xX
Ezn04kmEcF7eWzTzFI4McEt1lGr3ph+XA4WN8Ia3v5el096VkBGZSU5x3e0z2X8z5TxmoiCDirNi
NdDSiYVm8je9r436irfhH5Em8N0RBQNS1d68ZYc9W6ZK2Sn5WJa+3MJuntbzMDkE3iFQapOLAAsP
lk5erQxlkZCtoNKULbpw7D6KRuacAcg5BaZCjwHm7aeZmJzj38Fur0uY6Sno31xpJ1BKwwA6wgw8
Cr2QvtHzsQ3/yvaNadwCwkxpqUHepwIvB3dU0G40trgRtZyM64lsdSxtpLznSJNqLkg/HdAtReuL
be/xAA54vFjrRypLOZvE4H2WVHUmo7Oy2dT0NE3lWSslMNUKz0N+rpIKdQiaBEnop9InIYyEHMWC
hHTr81Me/FoLUe7cB5rJbP9hHfP5yo+h3OTrRMv8dXh5Ef0/8RuK8SbmSBd+wRV5FNSC1jiy8Y8W
aWzUMTubxkRE+Y53m7YKKl1jRjXSu9EYa8sRc53WGbtYepRMvLNnx/E5JeC717khx75ugfO14sn6
yyMYTGM4YJFTFGwkKPWhT9nirlYtR1AUi3FolpBD9/QaaqR37vPThY2gYe7IgHOWYHrTpSdKT1Q7
E69yXNdK1cFee+3JgaLUOVRoIVHZ0b5uoviqQPY6g76mD7Adx4XqKkDU+ebYY2mr0n4lmGJcb1Wj
BP6JV4QbyBZmgUfhb/ySKNnqBEtz6IQ7LczbXlMlu7s08pU+hIDTSbL+kEKTKPm6hAXbU8X12cp+
1hClPAdzM28cseYX/HSGp6YVwh23iCrLEMH6y/anirPgqUAlL8A96BcCKS2Jljq86kr8AnImfj7R
MvYwOZngLPXF4pBzEuO86f4ugVl0XO5uPh35b082PJttIh1jiaG8C0FGJTnVwdpG0J+9t4Eb09El
jMtVGWL1U/zNpoG9n3mp5qPFvrSUUEv65mCOqE1obKMEfRCpPtV5wvROZ0uEfvwj3kJBg9Sice0f
HHCLDxg/AvAnLoQ5OecRiTF0tQIDDhmy7nDpNYBDMx26YyqbUOpKneSOPzNr4XBMY4+tI9c3GjFf
dsL/cLmwDvF4r5o/2HIzrbfasnW9G7rbUeWX0Zu9wIOgtajPBi5g7UPHrvUX9QtThKbeZ7nbN0Ly
RwqP4wpJsELOeUWR8sV14NS2C0R5LtzFlrBOadAOC1OtZh51kLcwBIbivB7SePRXRSpLBLMg3TO/
bV9mCf3jk/JwouZk0+gajQihFv8P46Mi9EfP/6fb1ZEW3/YNuWrO4HDjnKEpyOe/U5jILcd6Ea8Z
jm1yci0SedJZJ1SxZ8UPz73zmnrsQIZdzIxkNLaPxxEV/nD/TOqWM43BZs+iebuJjtoutuRMY0Rn
ZfPWBv+DUZD0MY2u54YRBurrMau4dZtf+P8qtRu6oKyL4hXfbRA5hWRhtPty46/f6wJrMajHBdaW
R2Np80mwOCnBkWw+M7ifIoSU2KEip9yuzQr1L/7iu1lIkDb8ezhln+GJ9AqgbvgvUZRU9TFy0vjl
cXOsoXUIhIGiiNkhA8ECVoj3BBiWx3UHFwH0CxDWni1SP34khlHfAAk4Dy5KX3nV9u6acr+X67x8
8wfRvTjPNj6JXuvAThNCn0r4GgCkMEYv9+uPQuHBpWNODn8R/xz/a+P4izfAT3fbMZkSWPuCZlwX
mvIoZCzB5y5dGQo2X0R5R9itvhcK5pmFvR8mQ3h9GQ7BA4eFlqAnaRxGbnG8r5aOYndmSKt//iSl
ggDNaTNdpMfZTqibHVzvxBUeRv8Y3bLZeIHkY6Iur8ZGPM3mX/exqPD6V373sWz1PuCoga1ANdAo
3yTRao4oLeCUEaOee8vaHMtyp27mpogn9/lRivxVozWfGPegulrZrUsNa6YVQ4j+CJ1zeHXCZ0CF
LtaxOc9Bkof7vo4PaAJEWqZCYCwpnXVSA4HiTbA461rmudbXItug2Rvomflsud8NPGiaNpMmE9xr
qJzLEn6e4gX1hVu9B4paENzG6Le38NPC/qDWYZRSjDC/brxUa9FvjLVKkwe5svF9v26mDNX2I5u+
l8DgTjRg9yqkNXiH0PyGbGke3gZh79+X684/+IOon0OmNp8ALCTZifrYlevFtnNlzlTUVRMn8TNi
P7QmE3E1N1alqc+kDsCSaY6IFzMTSjqJ6t94x9tpsBy3PNvtglrP6LIHaMZouY3uMfuqQalcoUl8
UBGPXuGq/6y6ko/+GcPRuDI+aOTocSrZgJ4baseK4r4UGrNu49Aq1jvjgPHVkyR2J0j8/R5taXim
viz6AobIfbDQQDCFXz77J2hURpF325W5ouhTOtZ84z4ZUxBqjxHN00frz9ddoS5DyZia9HK86NxD
RDAEzPVbUPM/oUwc1YD5ec1HzXiRwPhcsyvBsEFOAeDnjz7lIkucdggC/snjcx84l3b1edjzrc0w
unpFQC7z7FG7mLUvq6NYokhqQORlQ7SaC5LJs1PvM+NCvWdXC9CIOuRhc2xj+yIpNb1VLNnPR08A
SOlqRw7bLcO85IgV7E2jcsqgyzumTx9vxYndiMRK7o7LZDbM7ODQBdHHh7Vov4wgLHjWsjwqPY/Y
s7/ILlseEe4Yl0hTpji4rs2S4lLb+g74X/RZBcE3JE5bQQCZgY6dXxAahFQr8ds36HA91c9LL4u/
6OznA0kjKHxF2LkR2bu0SL20KYEiNRb+EC/HyIuIJkLNbS4o3dYN5YS18reXwY3HW9eVhIjimo9D
f7mF2F3dByucrik2lolL/OUUR7Z/kpSswYvt3DqzWZiGnwGyd5LEYdD0CEIOw4zfqsZO+oKn/U85
ZXhiT3mFqd75vaBLJ+13iyF+ZeQip5Dsw35CebzIv/8uPaxebpScD6ookJ02bOVxfMLHXjCoTeGS
k7p70QCkSUojIxj6I0pPc3zxoYfWy3mYZEUzeK4No4dVLEIb2LBTAKVtHiasDdzVzpvno132R9ZX
oXb033sfgf9mOdlWnBYagLRMJHRP7teqE9jgErRE9Ckmtu3RdXDHcDHaXoi5POI602guzVg20PnX
FELZ5NNPADA827q10oibpBWlRxKTvxfDpwy9H8DnhIcM+3NG6XGSabRSyX+jfskTlu8bnkMkAuUK
n0x0N2kE/21ltLiV6e4dt1K0XJthEIf/09UK/po2dyAnbvo8Oc2PfcD6LFBjudB3jYWvqqYn9ozN
qtqKpq30QaHbj4H8GXzM0wLESRaQ/A7fk4+rn32AZfhlRLK15De/rTZ8PX2ON36XPJdyUfcnktu/
pu/SSr18BO4rrvNLBOQ9M6bmh3Y5xT+Yt7HQTGVTJpfP3rGpHuMAWfoKVGCO9e3wbFfhMLVe53Lg
VEu+HNoouYF9AwZD1qli7NvKpq4RQEhjvNFDvirjt1mGrNDrmueBhfBneBt/WbUy7QVmbDoZPuDE
lNlhkcKJoI0TQisuJ9ZHsBkJM+5DBlSE799y2lT9c/aOk40I1dAGGDuLBAxS/k/XKhS5lb/iw+ht
f9fZlPOIOdeD7tKo7aUi06pP8B6pjjyGZ3Np+nFCtUXBBibZpnSMMVxXS46SEXkAZ7JhpNsb1OvB
ZcezMNyKmjPcH3eBiZi/BNvpK6svtQwgl9RIqGKHk5jdlevZVTbpVuSa9y/jE2AVNLvGbcs8WqNe
uQqc9enXEc8/RmqH9pc4NZP3u79xayDAFLoeaL43uY11gBPc846kk7+wsWZswxcZPXBDlgNi0k5u
BsjETf7aw2Tdd8C1/0pcj38DOqAVve+QFzmpduSk/GiFa4zf/LHt4YIxtdoLjNckxnV310DsRI5H
38lcKnzWtxukC5TPvmft1OKpZe19fKC9AJKTzX3+AZP1aKHmViFuW9xMRjOnRPoMmMLaTxmIvZVE
wLESgx/vJUryDxN+MtUwjeNOH7Vag1osSwYFguQSzyFiNU7jw8G8ITU0N5spqK2hI8jrVs1Y8RrI
2J07FoA3bgs4gyHnZ5MeuIIwCqNc+OVhVAq+xA1TDzMrQfR2mLOWyzTWeWAkH5Hm3RR/FkdioJu5
fSfKx+iPuuYIhSOrijeC+m5F+YNqcTaFPAquJGsRUQFeR45NpifbhdLPG1aoLTO5w3Ouy8ZvuVqV
l2u3BO0gVkJXzzQ+rK115bHZZxKoXoYoSQdyXEcv8JpJD6S/ypSikk7NmJNtTflLMwKMEUOZtXpU
ike2jafOI29N8NxU6Olp6teV8uEdEl1DawIKH8/dnjl3ksyuOHdzSmc9wobg9uxi4JFSzTjtJ2RO
qjNoN1N8QuUXowiraxxLNtHMnoDUOlP1ZrUgHSiID7ahMt+wdZdt0Th/utrcsR8qkTOHtl7OBlMa
OpMWCcTYUk2oBfSjDMWp96JfL5885Qzfn/9Vz9feSutsYX7H6jL3rIdxgWjsiUgTCZM+ZmqI46UJ
FEZdoaSllTOZ6Z8gw/NpKG1V53CW2PAoQrh6R7z6Sysb5Fe95PtJemUAxMmlzDB/gm1PJAHMkwtG
TMOE70jbAyOiLvANh6pYquDiGn+O14uBH4OxsCveIOOkchLQouA8uamM7obndPBXFoUp3EI2cNC3
WjB5Nnf0rEblSf1poUWfgOoMrJq3i6opZyxQgbbAQU4/SgbDozX6KKRDHxBrJdOEO97bOnrIQnUI
FC5zOxQzRrlewsNtO2o17kcr82IDduUPbURZtnriwH4B42P3up+XoaoT06zdWPVv/SkwLxgCJn52
EVwr4L/FOb9NSEbcBo7sFJjRTKvDlAWIynAN5q4VJgU6UP7axn5ToZubJc6GgEqg3RA9vVE6xiVC
w2umX8PtPPXWfbK2iRiJ+u7YOqrltq5BrbIJAOMeOhxGOhfryC8zlHnJcRHiOTynEPhBxbU+6o0O
4xU7WWKJApVaPkaeLoCXNaKeNIxbsldME9M+Wm8Anz5ho3TK7XIhap9awaFSlFl5KVNyKFfhOVzi
Wkbm9jtoVBWWI3cbyR2dob0zdNH9+d3BZCVxuspVTBKYyPLxGR/LnwylnF8Wu4luMkBHOtZsd+CV
vPWwrtU5zj3aeY7vZlp7oFevzyF9pZ6Gs5eTPVw6foiqPtkE78+cjnyvmqJxhKDtpZVNK7ZPnNxc
zWwfWafwLBg+IxZPgIUscI4/+LSCFo9F9AOxA9rVHsS6VUPtxLmYc33kbXtKOSoOh6wbaQexZb4f
musQq60DZJv56yBZvAguwln6WfIV5fNniS2txqTHo3kYGUUYJDVJU3oFz6RdrEeDQGaubTVCRP/3
+UZyr4Dej4VYkDzc6gTWATaDfyz4nAq8tKL1fdKe48mh0c5oEdbXyzG9lXNQUNxkDNYO0Wpn/kDs
5tXg7Ld+lpcpSsj+sD8tAzGIuGgPi7TNQc5j99bPlSpACErK/LvI3Q4fT3sLjN3WYuXJH0y9bjJC
RUOWKAEuzf/xBB2ZgwyHomQLhIbFkrtHYFFXyNIdf9oxoRldmGeLZ3c/ufxq99x+GL3jJ1B1QinR
Mutad5Wy1dXcfpvXiEErbH+TUQBxC3FhLyWwyjMUQHhDLgv8VrS4DkBVvtK7X1Hm5ttXzmNpMW2n
6fpuxQVYu0EVhnhthIeDzRj/NwMY3tGxnoN/bBhhsEmYvMO+/25rerRjOMdlwylPkHYldKorjBqS
OoXuVxuVpCYPrGbBH40LzfJI1bWdUg73HoN9ZA+d+DZ0cJae4gln4J4RrDj+/Xf184I3kwiRmf6e
UZkKRTRZQxnO8KUA0JXmgUqMd1HRK3aRWDUswgvIg2fsm/6HHkdJSXvr8stojHbEtp8hB579HwTy
UgISjsWWeMzetLM5S3tYM5rMkW3XpBwtU8PWHClGh1pgtAUlRb5Y6myTXFaOr0xFqH6AvYOlyJwu
WzZA7LRsvwe7VaOFUpHMSO9MEFIJLcsRYC5cCZcjoYz6Uy0DraJWGdr2CTGrBspXA161sS6xnkzc
T5LTxY9d3ErarUP1xzh0t7ccXc0GajSgnchl/J99ggM8Mt73jqZp5MNEYfiu0hVxi5kcpkFNtdm6
a3QCj0D5xAV/8/EYs0sRBXasjsAOVpY9B6g5nsOiVUAT+57QrgBRyzV/VL6mX5/ZUkkhTv3ZVCr0
cPw8pVi6AOzHIJ1J8OQBRmFZNerL0T1RoFqsoX4lZ76CWsn6JVHuiaeTVwEi8YddgQau/dXRBcFc
PbU+DRQeYUCr7PE+p+84w9xWSQm9OT6PN6JqIH9kot/xLRsQWfko5zlx7CjgkZHIRxJ1YQ81AY7f
q4a+3+rB8u36A6dEjmET1RJT4WNMmyvltD99PfXTTfFhdrMuspuUV69V19ihE4PNVMTjjjMfGnqK
tb6J89F2k8eoW/3mVFKhVgSzbkJXfSAwsQUr8qED0FdwfYj+QbgYeOmC0wY2UArbE7MvnS71SRKN
dfEqmUPOsBAqlaBdI/Sg/OjSebaRmzPw8SWgWsLyvZRmeO6mAk3ZGXKuy6MsoJXnpIwJMwvHI8WP
b9O+RtbvfPpQyziPce8SCoLlfBZzrBqoF3wpW5gKgCOqGikFoip2HNxkPrPZa9t5kjoGFjgQ6U/A
1IbYHpDRLvVXGdxsCk9drbzD3jtMj7v/55trXFeHIuDA6++xysxz6FO2T6D1caHHCZoHl6zS7V2v
kO8inEKhUczmzBzXCz4B2HqYV/paW6WRiMkew9MSZ52u7npiO34piRK1a9/vKds2pd8rzIVLOQC7
VfaskSERRc8EvpJAG0lh7OWxSXu0HWdNB3gbL/MNemNC7VrVsuplm6gqNsRRfm1qvxuYjEDxt6y6
4ABqp/KW3rBnxXTYu9OYsb343+045PvDUfJORyqmlHm6sbrfB417W0ZEJ8apjGSybcqSiZCDE5eJ
/bCi0wAxkWL618yzobKA6uGCO6xcHq9/W0k/mUzDt8s+YXzuVwi21NxwlbQGvpcYutIiY+vGYNIN
EaNtAiQwlqhBJU4ak6Wz5IPBX49+4CkooWwxR3c9SOKAVBXbf/FrS+8M7BVZ2p7wGUPD8jY/hXMu
gUYo3k2YuE/Za1KJgohxEvssfjBcwOWlEg/lXEZ/6hy6PnP693q4mIs5jSBkAanapcYHeqf1IlIk
d2w/phUMTsR78vdQthkrOgUvhwzkCSN4jK68cNF2vIrhADNZBB9v5i8xxrYpVRjpfBsf1GOifmU/
eSVq/TNIl6k2N1sV/h31eakt7tIesDos2Top4nm7GC1Uz4VJ6ZZLHo90gj4gpkF+dyjQx1w/28Lc
/7Hf9A6ieydpUf4JhReM2wmZPbWHFDh6+NI9Xw1DuAL/xLUt8gCxJfYo4nhQ+pxqPWXHg7yoV20/
L6OeMbTN6AVBjfANNsqmPMfbZKh15g3nvPvObEwAzuaxyzkuG/bJOOUxlz/z/XkoKV1ibTqwuMq6
0OA9ibtevMvaIZXBRD7LyP8w0JW+949b/utpzoqt/l+eZLyE4fXPEGoCeZ9n2HMK1tUTNar0UFjD
d1KGb0XOkBns4vHQz5INYGJiMl/fxm0wtaeG6L/Abv5Q+QVtEH+oprp421i1sMULJIwM69cZdR8/
D8VNK/Wih41X0TzDvvx/zpAeWXAQYrdJ+JzJWBvXxrp7RnoTGbAX2+4uQk0/1TjWRjseKdSChtuO
QxKVVoPQCpkCUHMp7355yG7U+8E9wr34A0TTmOoMvUGpKNTzV7gvgXSb0Tah+IkiiJm2LBR0uIJJ
Vi+lhOM0cDfFRFj0TwrM6E6z+VcP/JXJB+IO/bgXgsdCUd3EzijbC+z4TTeauJjzxrRNkzK8NTJh
tsZHo25h9zqPxnZW+VF6CGto4yu1eh7Wz1wK7CoCxtoyYC8+T8mWNPCjY0hW09WfZcVUsIWbNTUD
hSmR9Xd06UsHjSI2psviRlxjgLY6HzNxe0evKrGBBNqTbYIHcz4sVN5g/xWBLxspHLQMi/jK1LSz
Stu0riGK9t3rOO8xVnTiNyRrcwAhgTJp5IcoEGdKmgrVPPgyFV/GgNYYhjYLWjiIPUIg/L5xN3yc
9xXhrjybmoaWwqjh8c0CezWWVOPsGBlsI8iPKXErrw1ZNwudcPSXyK9oj5lNQ/0QUE3o9CFVEMTo
9yNe56Ywsnau1s+NIsX4TYTT1TKbHRVciwwkMKtexfiqS6L7HbfCOcgLPuNHkZ9JsOFQu1B5fdux
mfhGbQr85obZVeUngNAnfEGs2PQwSPbRA9CAdE3edugvKxeOcRcvtbzOLwkejcOBGRrjzvUDbJd/
T3KacsQhRX2O3kU9FivvYvXvdMFavTQ0z6scCKJozLGnRNuAvWLT2rGwET9l08kc6KEOsolDbLD9
x7WHBxVnO4DLUbn6RX/HfjlNEwEfD+yWwk57ZHwAct70NPnfksdiQAi4+bjwVqA7x8RdTP0kzWg3
04Eo9EOlEBXaG3F9ydzLYYNa+zRjYEtsda0+yohl908hNCZWqMfDSW1i2CERNVjwkF/on4FcHajy
RmpnSHzm53H0H0V7Cqi8Dij3R91bo16CoPYO03p++jOff+X7eYsT/DuyAAdgylJG+7n5fPuIIlpr
tZPdHctsj4A9Fze6Ncb+LmdC1B9rMqMqHnEp2QwsEefbxpHfmiXj+i5j8oynfOhc6l19gscVWuiY
MZn/HnaVZy9m1/PMnjqMs6bUyRbUl6BrpTtwIZlnHWf8mXSTei3d7+It4wLimflJ96Zyw8Dw4/RT
6gCmTyXNpF0vBd5qGejk0tDozx6N0tdhvob5ZpDyqkAmhldTg96JaF1CT8L5Q4dYJVt2npPuOSJx
Lmd2kfsk9aiLYfvgzphKnwNBnTXoRM38NoFMVsj5BlJwmaAgAATe/fYfDNEOtWBMuYITFT9zPDMT
WPM0YLbdiaQVw8zujlOORT6mRXfgWCJ6bTBKjCh4Gdd45hy0t08Hfg84msuKDJmOgpCR+UWvs0Ja
NrseK3UhFdR+Q78eSbDR4QmlsOMbDE9b+ysuuaNDnUJzt7AiJK7cPIOcui7VMyjOJpL3BEspuY5w
thWTD7q4XzI2MZyh1bbu3LSAJ4pTICbgpaTJwUEVwtrq9ezigkmLlgQqboveDqedyeHatwQAkvPu
YdRcFkfGu+gWxacFYmTd/bd4lzQobGrjnpjUZwP3dUBkDoQwlU2XpcRallJ+aGAw4y9FguKAXxZ5
dyfmvO4vDFshplZYfw6sp0Qq2PZeiiJUJvBS9efwpnDk8Sn7LpkdiXIOSBUpxTsLwZL6E8hdEHH2
skfg9slojFhXz4+rccj7wie0thPjHhdHnvyDVHadSMUIS9zC0FORMbdcTJjSGi3/PcB2WeVhPmHT
C0iwQt2UGF3yl7n8LmuDd6HBjJSvZN5yUNSvSK4ileGE4rkhd2y4HD/jHrHQqTuJomWG8R+zfd0O
GdVgxUubGQoDprF+JWqCCOKvKC49et/BAggH/0OBvHGHi1bFa3HWThZ8yVlMrOHEyiCButlMMoBs
xxNyjdpwy44+gh6H2hkJf9DB7PMghuCN86M92/gY7mtHHPyi0LEj4KAV0mfr/ZQwA3y70PPUos35
RGKmtUpvQGBTox1soDze8iYt3RdDewHxWwAiFNfhrISfdH9mWi8DEfmDMU+GlDO/lgxi+KjryA6a
gPDAn8fyJ0+OqDeqd+lqWYHbEJG7XAaeUVPvmjKo333GxBWIDwdImNozYw2RNvWT6PY+14qhUAV4
NB+ECIuEvX+ugSq4TVuSduH7OpZLlddWSCH7SKYhWSljly0mJrasuSNEPSg0uYYJwCLOIggXdCbm
mPo2KpLBaOgiPe5Vq7XhilcZFVW+jAKxdUZKvrLfQn6xXvIAq+U8pTy2D81smP/wjR4dpKFu6G1o
gtXQSpxLY302K33tW0Ztz4Mm1a7fNs+Yvh/aBiw46j/U48Ah1b0wlmxIj5Ilfzq22T3Tgo2c2YQS
uQVE0ODnDTbu4VCfkoOd7qNKQmW1Sp5+QewWgCqtxeHcbynHp8E3WcYFqKS1hGFnXpEHAIAhkrUr
nUHZdRk6ZreRQF37v8237XoOsYV3EsNLFUmTySIEmCKuWrRduAE3FGh1iDzAzxJcbzH/JQ84bf+X
/r7y8dMku60zEqrZP0uB4yicDduDkWEYvYF59pVAgCi8oIRu0PlyXG85E5Ax8xLLptJ0r1hULoPS
6dRa7IETp4JnM0drFoL/aJSZrpJnPDduhFJonPcv75UnLooGH4azhe/TK9/I2tibCMLVcBPza2tx
wIdabOY/h0z5b3w6yGlqCz0tZ5dtfYV/HqanHquSVkrUsZ4DTnzxhoZsFII9GdAl9mCICwoOAtUg
jS8kpSq+0uP7ZHzm9147XDhTdzLXLoNKFHd+xW1A7dmmzo6QwHjByI/Gm5cXOJG5btnRonSyh+Sq
+mz+KNCBqsMNR4gn4WqbDBz2xNc0l7/ARbFac/f8qMuEPhsxswdmhqlB3vA9BjtMXym3NOSDlHm9
8m99BAHooo+d6T/W5xMUrRki6hQJ8IoFc/ALrRRdhZbBOKFKuKxeLEoiVDtMgfde0Xj6hsMoxDE/
69mto8TT8r9y5uRHZOyFleBYNRfxZBIL6s4FpdIcxud6dfN/02npyl/HxNrIDjIrwz3gQRLKhIiT
O/zgL4c6FIwYxItofxyY4qiipw8S1WtvIlKeQSoNQ8e3azAlUoRV24wBF570vortu4BzgKe7V+73
UyNCfDDHTgbmd5HI3yFA/PsGyt45uqug7RQGDI/RiJY8el65a6+7/IKioCdGMiOF/1o5HFAB6cra
5v4iKaocEM0t8+7NtGGb3+g/fgJBxUknfPFh3taekFGdKuilJPpQtWqgsPO0jxYRiTocksE9WVbp
VjGB7tWZt8obJ8TYm7SclErI7TaWu46CGx5qr8syhEZsziphNoubF7k/rivenX8H0x62TxcOlbEH
3vAck9RaKwTBxrjSn/e991/LMSlQ6qdzYZuXZao1Oo0CoBXcjYNGolHMQ/H+y9k20PNrRx5hJ9JI
tNjNPr4tTd4H6Fyo3xBkyLmJr3iAZv7cUyZzGAHb0nzAZOiQbQn6za8qZGucInhWryi1bvCfzQ2K
QkSDX8br2rxezWvl2yQmPv5I0xu9iFRPqkybAD2NMGhiZBeciP2i20HWU2re5jYt7OtoBerPjnTB
CyOgcHlxVo7hMuRJm25ncWGvQEBC4Zwzr31XWTFvUBhaR/AtoaQzYNtx12NSSgFTNbpVjII6He9E
IOBZoznUEY/EoJvTMJ4fiQVplybrTgy3pVBwWsS/52am4ecZLy1gg8a93yOANpXuLd1xychmqmBh
OSfqoAiQDk426+pjSqI/YmgBUz9MsMIYWaO2iBC6WX2ePcrh3vualuxEud+Bgs6UD0g5swtq+RlE
xK8onXefmnmENWHxCjQmmtCw1t/RK1hGtajDotat5qcTCXufyT4yX5ybsjXNmErCYZjcFNSZGt3V
+92wzsit8PfiMfC6W5hJWs0KML4vZGdr3PgPHdQuvtpSSn6bVKXLVLyiWEOcy1NB97HvJC9Gps4A
+k0Ovt0eWCPS1fi+eZVF+lCjtpA4DzNnurjuZOv9ACWbjyt8pTZ7ZvfUVargQ0Prn/967zb5c5fs
eK3BRTkpmsU81GKRVNGoviPl3Ga/9OnaHXxRoqirZ/iguQG7RlsQsbFbQujw5HEeZ3WkB75yvogU
cZ1rAsFedExWtuTAYWnvY8qf9jOIyM97RGQedGKoBLwKL6PUJwKP8RcVekaMp6x7XUJe11tYmDCP
sJzyO1PlNEazfAIzk5edElE8QaqHT2rL7gVthh+/gpLPkQKU5E1tmyQ/Ct++yiJIe66YHwR+JEhK
1Mt+Zg0sRLtQ07DywJ0DaAQVOfG5VU/pcae+0+2WJAvwJJC4ZSyeBKpuepDnG3Tyy+rpZUAkYJIb
L1P3e5tlM97avGvWHOYp2jt92FAjvrPWB0NS0dFDRqYCzHTdTgrMUBSeXzJIRDqvRN+3dViEQ2bp
gLFn8T1Wa38jEbB00lizD1z+c96PzVw2RiOUtLGXSNcNjsQU3Yhb31lsxDL5Bzs2d0TtbPX4lbZW
s7wGl3E+fLCfPTHq+YjtUrp+yqrYekNS2kRZG4wqdgN601bDZ3dpgFnwhKnUMJcAPJmzoqsxqf//
QiwyyRN8GVxdF49mfhO1xoTkjds4+JJ1lIvAvAvGFYgoSGWmynEJmo2bgrHORmvTp/1dshb0+6bV
i5ZPCiyoy7dOusk+NgO5oNPoISlbeciMe31tu2g8egxLiPjPgf3S1GKFXDl3LKtXYeCXIKiG4YDP
iAF/BpVu76bajsj3s1VRQSv5t32R6FPolvlbkMyQOGpPPecmqK+BcBl5qmz597wFPlDr5m13AOeD
aQL0vHdoqhlEv4O03UkGxgCkmx2Uz4Vm86M+oNwYQ8x8rLK1Bg81X59HAFpfuNDMhdfzJIBOmmnE
C2Ua58h/zpvhRNuhN3KNMpH2Xfsx1SnwNjZjckZUWhq4IWpHxtHi0hSsez1qMQoINYRbm/Lmxk4V
qm0x1YVSzheCkGOjFq5aLCxCvn0FBBbCkxZ6rCmcU+nQXX1XiDHbNomfqSG6SO/GIMhcjYXNdK5z
ZbHBhy+4kk21ecHnXj8WJoJCp8A4TomRg87c8Y+NKuihrp//adOLDwxo+g4m3NmBeMxHqPjWCCPV
kVXBWzXgtsyb0t+cKInsfz9BpI06bKSPCd6lrQZJGAwX1qVOTLtLJqC+VYvYYM6wvB5XRtfhnfVT
+uRKpe/rTcW2sQwNreV0MwKjbSc6zmAygsblPbpo58CpYRIQaQDK2NNGr7hLT1KL+hV1cNsPAmCV
7jmiSywN7dIv7zRvBAn3GRCrNdYsQFZmnZDZsCm3k8QVfCa3HgYBOkD5YhbkKQbt/VA8e3sUmIo2
a09XSwPmjFZx/bJVxKoWRSLdF/x/o29PiUyIIBduRC8zDrxTU/EpczxMxe9EadQPi5lZMenBvYZo
qg1ji2XMPpIWk8Irt/HNVlph9f7lbDWmAHRkjhlEjVY725+mJUOESc1PpYSQXFRYqiqE588eN/AO
flzPfgGQ7pNEtYLtmAp8sGxL0rCZuWG19S40joCx11RDaGuwoHabC2Z8rmD0CiqOuRJg0u2pvTtc
EHHl6bENEFIl7oC7XaAq2rRsr3yCszKK8zhjiOETuvnpfI+uxgCYbLc4MOGKIovCwlAdok7uaHNb
/uQQVNaZ/zuIC3Hw9KLLjHGtKMnEFveF2Y5S4QLAl6vXlRlYJQHdNbL0YERUFCR2HOTy8LRN3WRw
c8YIwGNSFtxWgffZponh70T6IDVR7Db5EHwyfIl5TDTSVoPiJ5N+H8lUZ6AT0I22zv1JXGZHRi6G
6Hiar1Aow7ZsNQj9My2aFm4pSRTUPTR+krCVmNAKGg6fLfJhQuFgmAujvA6ghnqK4tOPaiyUvFkQ
gdhmYlhk1BedEfj38Ih9rF8iKgDlasudF/VlZ7QluxhJmKvPCm9IO+rhFUOp0Nsczeqx9zzkPYLL
GyUQKO3MpOtwJNEOVifMyTM0v2KgzkAVRO6JvwPUXAfZSwhmIH7j44/gxlQ7Ityv7ZIpGFV7zYz2
CtHWRVVlNEHydJbakMjnMluQ5HBBSXh+TuW0QGFCsT5FSZS4ZTrSvRhfcaHSuuu55tBPi8U4NT+A
uzx9CP4yW8NmZi+sJmcwPE4m/DcVWNCWmILqSO2nbNAgoKwFiVp1RqswOL2aL4ps6CwjxW5wn5kF
0jQlq5pZmy51Lu0BQ7AjCbPUnmRJZ4dYXKqfFzB2qxFSgzyd59KPEo1Iu0lfM8fpxVk4Jac7t5I+
9yUa7Tc4523G0jIRaj4Y9AVXrngN6g8518/RPdW6MH8bJOepu+jduShh7qUJOUoRsRY95w5DGZEF
mdNIT7V2OLIBdlNHjYyGW4NZYGSMQRy+somx5KKclxxWfOM4ZiQQEMj+lBK9nImH4n7+M+uXZLZV
ePVKZ4G7R/G7FqAgg9KfULVELomGyJ7a7ivfLc+pfofuAX1A9dSsSALFDbZD4DMwt++Vfmryavs6
Uhw7aK14jBOMYO6qB1+Ua8bA0y2i0TNkd9Nr1YdAgha8+MZa2cZ1SsLmpd8cvjZP/iqIJvWEMWBV
1gMzFhf+FLqeIPFEB0Hpa6D1hKjZG4xCpvzNZdxgpc3mYpvs0VP58nT6/orcuNqmCDMuMZM5r2fu
7vqyal9U29ixfmrj2BNl6q9ZpsMxn4xk1j5cTNFa4+oe1R6NilEf8TBGwFaptz8SwG7MWJtbGfmN
+cx59Jinmb/5dWu+0Q46GlB7fD5A/xnmNlnNtpp38eKRbDSe4QOp3qIoWgMVI2znNkFS4zPKezOi
F8Mgur6MFKlRbPEO28qBlSY1E6GEnYKlzAqUBj4PY1/uA/PB1QAwtX6lDlqt2dzrX0yjZpN0fq7a
ARaYC+Eo6qxjQyX5eVmy+QXLSjmXpxxhOEwCBmmMUvBE9M+ixNiAXz1XiCnmLKgZ2IH2si1jGPAj
7mshI2rq9S/gDYsZ5IfHW+3bB0nAd4yYsV6QyOE0n9WXpoftWV4nGJnHgCZr22VGj1HdingBQAN3
n9zCts6ptMk/V3VO5aOfLwlQ2rknw9bqeCesb5dZ7dfHLNcqV3DVnd134IQE8ibEUScsctlmYzu/
iijYWV4CDvITTIHa/mV1Jfz1zl53hI/4hfRVpkdtx++49RHOVMP+wuRT06JvgRZ1SGRALCO1zQlB
NJAcbmwYboeVZOza5o8nxRgRCSIqDrP/9q1iakU4H1E/f9huLlqdiA/MSTcT6iyeatxRcArMAril
jt5DymQ97UslU9my5+obMY6Vlar1EfcR8NeD8Pfh29EXn2sAxMIePKBCM1xaBxbiMmuMVHsoRJ0t
zhpEAj2h0kdldtxKchQ5xU5PmT7kjhLi6Lk/EefAmALuZezhw1BrdjrL7j+7zQkzNu6jgdaumT0+
ke/o7CxkdZbYE6fMew1r3SQI3TGow6UcdRlRxQ/MmJRaZwdy5nvT6/9BRa0J0fyRFtUI+APigYek
fNRu+UviR3MCuJRAM1dVn6hcAJ1aBqHsJ6Y2dMLnkSJkdmlDgpXJM9kL6j/DlCQCoCwieuYYHSx3
eTizKo7nvMMSJeE26gPpcwm9xK6Za2PAcec5dPMvmzyx/AtjDeU502aK4ryLkZ0wllJV4JPKFhpb
cti3PRv1ZU6X64vqX6seLdVfO17xeC/HI5FENnwG1kdUenKws0/Nk0nX1c/mH/SwMwPpfkOmHMoA
qRH3ZZgvPvgbMeE+/aHV6aq2IW5g/bovLQTb/zxg5DTyCd7YB/5zTUhbmkDqHXZO2VPNKaXanRri
izgNJXmFtHstSJqtnEv3gYb5sudYhRfx9s3GHlK9wgMNvT/EjJ1vwP/7NO9Yh9bCHxJfoLmCjLh0
5o78VGmR6O0EyxzwdtqaABZXAySg6g9NOjgxisfp6xr+9Sx2YM+uG/lGKs2IFtc8TL4HntM4aKPt
IGCXbYise0G+1gGKVDwQF8cbY8BawfDoThbT00Gdo6SwXZW5WErkF5oJK5wtPQ1xqNIMmeyaWfIv
BsjUHwYFHKmPpVhiSz7KhJZBLducspBKOR5CZaA+AgIdv+J6FkESfmvjkepl7GgrhCl9aUflDRVQ
a5momHWGfTkOIQqiWXpYxuE/xzNYOTbOxNuwtaTIeRTS/YSjM1mYFESQmR0NNyKmgO+WdnrrYdS+
4SAGAOTPbHCbynDsDbh087ESCv4Ch62lzLLV1nuU7no3UFiW2jt5gkrfE1N/CxPeC8HUIAczgFCf
qtHhaC6axDTmlWJODdYlCTJsw7avVzr018kYeUhWner7btSQ4tYW4izwOFIwPQyV00vfFCyTyGfG
aCUnfPrUEEepBky2ucs0sPKLoTs0x80fwBaVKNy/VAXB4gcnWG1PUCQFtpx4KlnDPnMSu0mV9VDV
RxOi5L3jO0OcFzByvt2CWd9ZoZN7gI5C5NCrJPLAKR4RKTSzrgIwJQ11TJoQt2MO1BtIYqqf3wds
XhDlp0O91z+HZ1V4/0y6iFU8Qdu5aH/iQ6BwjAIHVfJrqu2EbdGuUvUf9Jvf1VraAn5n4m+eZfmO
gXHffGIn//3xN9zbCOVrA7+rnP6aaN/93W86hH0R/jvaOD0IMmZxs3I+rsPnLajnUhcqrzidMdoc
STu5RWg/x4r+5FhgXXs+ltCnxaYZgPUAqbMnjkJUopjK70vvUoajMy9rkKU2v7Su41Tjx7DXjORH
rg9P4ZLS8csbw7MN6JZnQHGkBnFbHcHH6KrZwoqWHeQG+3QyORNFWJyD3ELm6KUAZCXNjd5pdyQh
VycpxrczJxvnd5lqdWVUXQDBsL00Sqn2LGzJj1+EkLJV8/utba5kNBoJ/SIeGtuEdkymdUjBYqfc
pBGyQqnH9d/vl9UnYSodM258ulhTciwT3jFVtIRZrUJt/psMVchggOEjwsBszSLcM/iEEh7i0A6y
gRXTn14sJ3ufT3dy9dTakSDCbImgAJpDkKpS55oX1gCSCA95+cVYz8ac0Q01LEJ6aWQcj2ufqSja
h+VO7yoOii4fN5LGUQrIt9D12Fge5zF0aNdFZG8WJH0KSCMYL8Crbq0UJTIcV65LD7clIt5Lwij/
U+j3ZKYqpERQjkUFmry6xH4EglgZ4XYoY9v/agmOIFvgYxaTbypV/4zoVZE3EftXmJsF0Cpmf5S8
I1wzNgMgaXvKzLMMikQxSa+iabhFBS+Ej6OE3FWC+fgES9SDyUcEDqQfe94F7UFKBBmz6OTto4F+
yMDd6etot2HKwsn822fwcLUgS2lizVgvngaiU6tNVn3/Y3skGy9jG5nFUJN3tQDxLMY+Ow/a//W9
FT9wnKFuInUDXBnbxziTGbISZ+VR16vEzIQIxPWq3/7oT9zEwXfVaJezZGFNqf6IGesqyktEq4bP
sp+1MGX+2vIihTL0OZ+2ZU885DnN8f9i1UipqLKVsgavxtFlgcU3/R7XWrSje3KZbF/UMN9yfRM8
Hn6nk3mVkee0EBj1MuJzB5rX0GIK7xIgF3hYnzHhnurL/52X3ynFDIqveB3dQF75lv68sx1BADoP
M8MlRYSrc2w92fI0MGrVGW1y4jp/JHSc/O2ubvgu3r3/L9Ato/Z9+qpJmum/5R16hTJe9ZER7Q/+
sqbdg6UxCt9lF9Dwog+Cs0ebJ0YOLwhKvPxaquFMOCafsXqDZFeozsP7C78mp7+OLu47oeXGv4I1
4R+p/LBrlWN1SSCY08qWgCkmUAmhLBOJlZv0/ah3P+Gd6pnYT+tcWwtKJKJujlhMpHdGYlpSr8EU
5Z1PWxqH+CwdUnFZtLDL862mDhm5TQ8AOqKr2m6QjHxpf48/eJzrsLeS1F/DMWL3uVMx0Ztn+zZW
fW3wtUYCrDuj3HicwnV5TNrjbK7TxW03R1296l8OzaisYhRHkAay/jQUey+ru2/cQ7mCfMpwC+Yu
9sPdMRG11dfqOs3I/Ct5ujN5cYOLizJJR7TTCG9CCq2UpOlnZZAeRe1PTvZnyIf43qPs8vM4dPVQ
lvyDHhzuddQHaM8/AyFf7XhIaUMF7VlnZZvP7AoPT7rqSqajcr3vj/TRZFDeLILRYpv6SZjPe1Cr
gd8Bo8kyEubTh0afyQm3IDRPZtAFHjfcgH4yhgXF9Yys+x2v4ER5GjnNAWStgtMBrTpEBpdoVchX
51tKmoTyMrStfakWTDX7iAh/D/t9Wa8XQuMKmgNS9c5GJq8BFdiUNaCtBuuNHNgjxJflyE3TCx+D
f90YmFNxKS6UB4r3W/oojXA+IG3OjnLPAebQRdjmVRfiv0LEIblBMd1l1rwcN46HxgcNl+kaEnXh
D2P/8BbWEIogm+u1Exyv8jHJhmun8INb4T01CX83yYxCfhUza+bTq8wanUXdfuOu17F9XbSS6QFg
9z2k569WQ3F9kbkXck1ahBdgmrkbJSyu6DbybeZVlO5sQawhMOv9jDgBSyj0saauI+VpwF/69HQf
hRDedOQjXTd/KN5n4OkcFnDGnaZDfpmNT+ku0AwROqa4hLm9m/hT8NkvpEJmAOmtCSFnuCsKX1sw
aHTdDqc789LuXBlOP2hjk1EVGN6jP0B0bK30PMTEwuK8s5142Yuhh8Ci4fQc8XXSQBRMv79oMD9Z
FHffHUbsWJpse+CceUQTKkMLqBUlmNpoGYkXMgJ2YhILhE0My2wA/87RvpRITshv8RzMI2sayfRf
TvRJus4HonmQIgq0zOylwJ23UpY9hHiDhm3xzOtbmdwCWDD0i1BKOA4go4hn8DD5LfuUQcGjjo1x
4Vsa10w++mSmJKx2b5O/4ajO++mgwkaZrbH7lxl/vGwY8fK9W3f3qS1N7HABRRZlSV5cCG/vBjo4
ifV0q99Fv84RHw/Tu2FCZeKKCAsuZcDTlcFiO+udFiyN8Dr3Lki1PMu77RTc16NahEX8Fs9CMgHG
EU7QPfa8nMcEtw0i1wRXPZ9HOI67ucGTlTfph/04HjWRfGJi4ZrQQLGTPzqQXDwrKK5dVWsSx7QQ
tRZaXtfaS3VjFoQBQv8+v7mX8Qh9t0pYA0MdcOWeEb0BsDmgE9XupmRSZoSKEam8Qln5i/6qthwB
4BHXCJB7kdpw06qXAYQR2QzE7Kip6D+Y8XZ26U9l5qVDh6YD3WbzLAZKfo0uWS4jVnOZ2KJCyORN
3hgU3VQ7rA22KTp39JNdUjf3/aRENh367gRRud16bNZE1fxoutxovUS8J3GcQHy3gZ3kCMetxBEI
hExrR5Z6wgQkVwVq4F8V5AOIrs0lUe4qgZE7gFJGPWzsftTt+QwKaK+6fBe5G3eUBfVhlthV9hDd
IW2OPl1CQcsDyoEbi9yjP2tHWpuYch9RnmVo/UBzKJflj2XIcgriBYMtoCNTutDWn2dfnx0wFyYQ
1AHhu82P7Otv0jtODrKQZtuT1Cj7EGTQg7GkswvM85fFv2yvNNS6/mRZoSECVcLowB4DYuiJHQEe
8Bzu/eY9PG+Of+ETGTsFngum1ebHJnJcurFB/r/RaIVHbTbT9YX+ApPYI4Z7NkfRaERIKM37X+A9
kCg2nO1zi0B93URcs2iuHWGcBSi94UnRLybdlC2RkhQXfYcELvI756BborE1f/Z+/PvGeylSKJFP
uLHPym+FO3ufots4S7eFZ7Q15mvPzYuogVMEt56YSEr513OVQ5yVhMz071JzYTN4fjbtSrSqJzJv
0piRyM/9yqIc6iCQHifwT192Px3f6T+cC0OxJgXWCOp9g/Xv8RC7Zi+iw1Fa3kOU+n3kjAIuYEFN
0rXkDej1tEbjV3cSO8YO41NsDAAlp2H8hMu4l0zUrzBGoTeaBbjb8RJ16qp20SGu85PJhlXAcTvq
S0TWhmQEzIx4TwpARWWX9M7wglNKcAxxSdsuyXRlxzYiTmhaC6yc21xE4L6Ouk5O4qghmT91J5Rw
iABDAsj5ks9zcKnlY+6kfgtUWkn0hUWr2OPmx0tOjjSkzJmEF0Gj+0VViZ4UN3keNKBf1cwpF9Kw
+vwYf6hCGpTIeF+yCUQzzMqK3AOb6/ngRPcvwIvrXg2G35ZaA84vnmc1jeQHceTCTmfznfiPt8un
k+zwHBFDvI84HapxTr4NHd7Ijx575FEdCyR+I/+QuBTpzothphK1q+2KzI7YQ5+hj5M1ayVSySzO
x4UouXLnyjPKMHbe5e4A2pV4Qdzp3VAC6j5GRiKdzP4MXcpMTjm3RDF4KQIj2WRnrRnv5YQ3B5Es
g+IwqECniKTRtD0GRn1zTouvYh8FMklN8HF1XRwLy3atikInu7oAUmqsPbhIugd+Ebf3acuC3oKS
NZfZa0q1czRdF1Y74w88IghQbmbVVeUmAsx/a2pjhYUUtAfn/nTR967VohiclBgABp4oITnv7j7a
4sS9OkzkWqBibr+52dByIMAm+3Wp7T9oCF0jP6MICbFYnjIn3oGz4PiLF1pmVITT6iitUeuase3t
k7PZckLUIt4a7nv5bwCLTc7fQ/PYpsELQmiiMmd0d+daixGe0gKwr8BYP6JFKIlGIRbCfQdBCz1w
JdfCs+nqa5DF9VqA7ysHxD02rAmpV19KVD5YKYu760zCN+8AsoI+KYmn3fXOvW4M1VkwVIIeXNwX
C1hAQutzki5HCS0Fp12xba8mjZ4iX+Kh+ka67J3DulbvLK7uLwwiNGViJF4EegZU2aeZAEUVe9Zv
1N7BqJE2kjdjE+PmQxsKP3lH8W2F9UCR9eP4M3uQT77nCSXVpW+MzGzgHJLDm8g3e/cNUza+hkdm
a+JIy9eH0AU1Pyn2JTa9hpCCcD7sIuocTyW/RUgma+UTkF5+JuqLV+Occ2xvdMEjDyn6NpY5EnZE
XyC47hBhBht4iZNN2wGhEfOSax/ONX9yI7VsID5ephfPEqMw8ftyLN4XHRygl5Vzuc7ZdCJEPL5I
zx/EHvBz2fyWHiR+acmBS0JBSvE2v5YABlwg5b+cjFlchi4oYNyiIBYmt2x5NFV+Jnd9SRW3Zp+C
RzcxtEq1L0hFdzLLdNYHlOkO88Ksg9UvD1QPQECdm06aa6Dw9drnWhH+Q3WDNBRgjKQvMk2xzXjh
fDJK9PVqSF4ZCH9l338XZkj01uFGHcYehzXxvxD5tPAvqFQz9eHZJ6zE4W0eHZfHIsAGYBXEPwp+
+Cb2gUISVn93LBk4ScQSkcHtOhW1buzfvFutD7vrOSkLXQDhZbQRfnbLnlvcTKcnVfQN6NXDmSpy
dx3GF7Vn+VOoQcnbrHHF4R5A2NCO/egnlbV3sVr97iOsWt80p5YxqqOGy9EDM0N+V1zxahrzJO+N
6KMDKz1nBgribPQWupfleWP+o3m0LinV8qjHfOjkJj+w+3iY/NNc5pyU2YNzZQqGvjEtSr07b3Sx
iLol3VFhzdVfS/5C41yQ/qxS4kY6b3wdavRsdg6Q/rXkc73Su2yXORN/hWbusUbCovKcXd8pn3Ib
sqp7VXdsoZfNZpsvM0nr7nMxw6n0T/opnx16cF3aiHn284JRpVk8XW2o/pTDzJZBHU3pPsVlDVO7
CzQ3kAYfo2TP21D1o/STV4+P1zDAJg6OQ2ayY48ag6NaLonJEocF2rR53LOf8wt03gTlWoy/YbYs
G5fcEsf1unijh+fdSHnP/I3nDU4JZfrXPfBx59nNq1XHceJ7BV6sr+HaseZd6k2KSRDgxKDLSJd5
t/mvyZxvQwY6aHbcsFCiPE/wp5cEDGFM8HIX3bPmG0NpcBpPTpAtfiTkeDARxxl8W0z+WM+krlE0
WdBxL+BMBTPufuG2f9bEf/7XxjZ3fN8SjZ8vIMcMqCUX/IopbyhRLPrZDUX1Y2+lIt7j8C0N6O4+
w9xY7pryo0dOGrnVxs1UfI6X+9wcMN/96ssou82hbQwQoNVgA3pDwkaA8evf4txc2N5grhMTbN4b
muGHtSVhi6P6FD7Yt492k6dgYiHjHQ35SNHnu360fI6F66GtVG6zE3mEaMtrysKAvChpNujGL726
zeYKeYXujNEn6yr5Gnp6d6fr8RgO+Arn4ynC6q3d/RrEDhntX57geBfYiifZ/wEm8gScomfZVTRo
7TpkjmwyL6JXPZCQeo8VQ1/Jx1xtTzRWUKRhzhAxhDLLumQ9J+4dqF47nGWJrxuSkTPiNfMse1Ix
O36o0bI/mHIRIb+zica2hR+dYS4pNOq5zTk8EG2yiiahLzokTqLIoSc43o4HbpBCmKrFDThYNYnR
+Bhv81f3bZofxE/6b83mwZA4FL8dY/o/txcXcKdkdMyvgprVFyIJNwMsC0FF4tnON7iyuM8WW02l
Qtg94A7UW1YsQnbf/+ljK1xUYlGPlWB7z7dAiu+T+xjXwYJFBh/6vKSe/fUQF8f616qUoK2dPbPh
UEPbUmlThmxASYuDU2FZZ/4foQn4h9C76yoWzNd1ANuAX41EcY7ecB1WVf3zugGRtY6ONrDdO5UY
iEdfmkOkWeqVYVb/9w9bglnOcl/gY9GlXj1qSfh6DXk58J4Ve7sebXfVdIF0JMuUgoRMyOVIAvkW
CYmoyJjck6LAfDLteGbMl79ktC9pVCZkcru2xgY+wFAYmp5iKSRFMbuwIRQaZNr2JgpIK+ngKgxl
cWCVt8Yq8rRuAZyZ2uQqP3WVneHzXR2MJN060Cs8xY4nTYXBjYiSoBVOsB1kQLi/AUpsQ6tRmYhW
ZcYl4S9nMjJDadbz3wRT1Q+V/Hg4HBRMUnzBctl3C/O1KqRaX3TYYPJ7cdeB45aRs8aAN8QB2Nzn
1vUOfAjHxnngwZ33OTLye9QqwVAA/y5yXC3Y5vDX+n4tdwLh4fXuzgcW3CPvY8y+6/FnuqT/7JAl
C1fYZ9yNkBxxHWsdvSYJrRzKB8eQGBDvDJ5nqcBfhdZnO6m6RgPvDW0kY4gUN5AGDdQqcBrhID27
W5UnEPsdsuYe2gsjmY2kLXaAJoUHJHTkHUDj8ZUivLk9Jlwd3SOhpeJKqrePlWulgxydL4O3RD1x
s93kZlZXHQRE58CrjJ0z5pTtfDmlOnHQ+DhM3pZmRQhIpk+qvdVIp/aA5pqRWQg+VlCioMW3gVSU
1ROJRpP8ZQotYrwa+lsDskAB6uT/rr/KPC5AZPc9YaBAFvUMmh78OQTl3LGffb+rqrfj65OTCLSH
kPB4zUmTFmMIrmzHJKYb9hwZ8G0RIHSPegqEbyth7dyhp4vOS3huR2GdyTd5VnEKrYKUNo7fysQd
54/KrvYwmfS5elVedZsymQfgIunlm3mgsDBb/Bj0IFCrqskLUGKWSVXQC5PgjMQIvJ4kc5ZwS5+6
YC8B4/O3K8rUUpkDso/5ou4kayoo0uj23ANzXI7tOYiPf7E3fDNROMWh46Nyk206bTgzpJU94ziT
HrfTiS2RgL1Y8UKWaxeG7TJa3Xl9FECqCSln/HvcwRLuBX0TxzW+3XYVAeqztTSCGPzkTnf/g+Co
1zObUznkJGdvIsELHXJrzaMq2fEcSE0fcEs8JfDYJ53nKD7Uy9QBhmh4xKyQUnoE1Fy7S75gABoT
cJVO41Lt84503wD1bdpLLmgkY16pWydwfvLFvcTlTa7NfJmAtXbgaQMQpoxX2+PPajFi6lpj2Ddc
WAUrx8X+qeat8rFgk+dvgV6BGTZ8PDSho6kaRyt5zRh5kZWc4rPnBhB3RMES95bypa92hBhn2yO9
2u8IgKhiWsMj+mHSt9pIeMl0tTPZb6rATxtx1h8SzxvNQNsoIhb4ZLYoy1IX7t0J62eAlNfYx4MS
NBGbFpGlnD+B7g/odYOYPvc1ix/p7IXkRimB51glxzfw4fA5MTpkcG5fGSepblk9d+TV0th00tI1
V6tUvb/gk+8J3ZXGhi5u4BzLNim+0Yq4AE9CqJErKm9UIg0KoVVYpWYWiCsJY39eCe/dOYnpPRyR
vBmWiHHz/xWFIWpqWJRpzlAH16Z1btktRqik0NgkzimwQATNHh59a7FK62oSbSlMo+u59rfe9RQi
IQB0q0gtYCBm1HpICXyVjB0FBJtQls7cfYiDng56UJHdkKsFQRyNJWftjwVAaesgdP/PIUpd2yXM
ZNc4q7/+A2vci2PUY9a5meN6tFDSS0G0J71aKCh2rRLrs69nvT1510m+Sh9bekl4P0VHBoCfeYCz
cHvfSiyC8NFsE9olbHwS3h2yXRGreLpqzW3VCnSEfBv1YmZvD/B/f9NwtQfSZl3BGopPFi6bPT4f
/VBQPaQHj8j+flfIVAdswD/asuThlByYoedhiGtqRUpnc9tFaEAe7u3PGsj415DndzGVNQTNCjL3
IZeYm9pV94zYpkCxLvRv1lxQMFONIw2t365TnF9OTxrxLBkiNoImImz+SsBZfX6Lbs+8vdrXBv3B
DK5wfioenkr+pV25B/hzCPGP6HLL1wKVTz55yDXFGA5suXtvVTsd8jx61enq8euoMGu6yMRv/Dba
/BwhFQaPI7EzapVdaVrlCGsukznX3ilmgNK5hOR29e15Jdk4vaI3ELCW9ZJkQWkL4a/tpkSsx8h8
GTBEx/oP9QC8t+kzi2xbpbFoiviDhmWVHFSiJJW2J6G3JMYOE29jtI6QOfNs0cdytMwKOdDTBSri
ewlSNt+K3GgyPNfyj2pWUxGBeb8T7Dw2DtD94sLSFMxgsr7yhLcgDPyBLLN/TT9yGnXYcuBqDhLj
RJDqoroo+fPJJ6EDfCZKGoYfb5aByB0SDkDDigMNyPDghmOjTAJXLriRMPjoDd+rm0vW3I85rNiR
YeCUBn2F+8BtXOcgKKwM6/NER3Y57ahJrHUBzqVbM0RcO7xAttTTn05yZGd+shU+AjiVsMfezadm
/n3GdjaUmvdn3M3sCoa1OhDL+yzfVgvH2lt9ovUEVdVoLV3fENG6F7objN95hN6Ew+WJmeJ3wDGl
pMzae4kH09JF+uuVFR/ZE9NziDfiZUsGENGXwrLgxf3amRLBNYkOAGAQfnasiUrDsE7u0feRCyIy
liAbWT+AkTkEsPSHRk1kqKlZHUM/RCaaDi5HnVvK64k0elE0k+bpuf21r4YtIYmAXBvS3p1oFuOn
wSiRdCHtoRG8czT2YGuwehhpGQTVcSsGuLeLQ02u3/beH+eRS/tkoZ1ORSizh5thygsY3grcHym4
JHUktScFe7rhj3wXEo+kjyy+y9NeddtwC/vuMz2dp2V5C3TtpGfrqOURvcKHGjdib2191/3sLKcz
ovbns3qVQm3TRQhtZFjC5/V3AOVI6eazLX/r80wkHIdfsuuthz1WrOl15ECJXs9MI2VN7URfOEJF
UPzvFkTks0SHb1RpAJ7kLwG+AjLg59Zp88hYzNtnfYEAoS+PDcaCBMrqRp4MWOAyWtynPl2Y9iMa
QmNKrUdGs2S3qWRwNVVRxM9gNeJFlqDPyPlgZfKTPOli5YNCFw+kzgmuoADuAzVnHxXlRXak/K6g
N2QwRGW2zJy1RoOHv3QMSja4wsiqVA7UvdE/DlDg2s9BprL+NAzeuPBFjmL21mjmD/KPc1RCg0wI
P8Us1pNyBadU8/y6GxPzIdgw3aLYU4+zEeH6/R3TV/F35LrFeCqQD1JZ89SbH3wjluIY8j6ufVX9
T5LJbnfR7KKg/tWSEkJWiJRm+7I/mm6+VmbG24ytZVIjKCpw/YRWVtdLUcuMZdDBwUJm7ovMBhds
vSpsdwPsESU+yrw+S+dOgSLc1I8uoWGuEkh62Ropls25eInq5BbRer1Im9YfgVsJJADYpvlZViF2
CXbUcVRZ3Y/1RZZtmXUd/FQdbXAUOfc32n5GhYl7zs6K7wJL5mbkmSuweReUFl3WNfv9zLkQohlB
ADco5mnGfwU6FhHXmo1tv9GiflJQUme6718WBQfAgCshZgGdp/tF9votZyVfDsOvbksoQZ+pGUcZ
ek2yWd/PkN0jHBsc7vNJMm75myekTdlSPsIhirQ1SQ+RDsdS83az8RyOqk0maAS7LV/oPUCNSuE+
nGFK+yVR2ikmIBnQvhDQXDINqTmxkcbiSkSCjCEAGSzc058H0iablUv5dJ3HeVQyZyQHnv0vOWdc
SlX2/+MXtUOnxHnsfhWBF6eSxZAsH45kS80c8TGDJXlTUiBACWY3XN5yHLz+RtMMwPVsSV/98v4g
918+u8+4R1Tp4S4oiekdE0KzIv5PIMDQEyYh0ivSLmbSUlwFqIH0OHzxEFu+hOEJB52aBpYxygF/
jxt4qjXFVeItRpnCyBi+M5Z7odP/9O26BK85DaeuhNM8vXE52xoPO3rM2qee/DvCOHBMPagpAUxY
BMnKkVdwWQPhONEE6OlcDBrsZyI7l1I7oseqECZ1Go8SkhpS0f+nea9APhgIjUVh4XqAyZEEEDNn
SbFnyygFXD43CB+wxnENHVsG7k5PnhsriuDX7mRB+XvCBPHHTPiMTCSauOzMGOvroNgIYH1eK1OG
rvbbZGxkgGqqSafMfwshjqvh7tD2o8OKDH4ZGGXMTJVRSX+kuBHrIDZBEHm+8Z/aXPchd25eQjC+
DdVuWxp9NJx516hq+wdYC12MdK0OFtQN7f4VYJE/p1Bs4ceXDZgCdoT+iOOD293oLg8+ga8bXJ4B
Sk9Tj4P+YshVngrq7+f5/U64PhAeePwBTPm2OvLiR7rhdAEvkuvjgLTZ0qGe5iNK4jNpubcWWKvK
5C6Ag1EGJTDI0nwDGiBtyVzRCe9DD9bJUaEPO+uX26QeNMDSzxR7ejfjZn4d6VnDV8Ban1DXxwLz
XOh5XWb8mBQ/ug/44eR1TV02afMdc/zKywF4OykafzR5oUQ+Xrhp3NPEj416ci23pTJeKT/yQaZF
KG77wSAXkbRUGmZEiMv1Kf0krwgac13rwu2q0NT6ep7DXHxcAv6d+ZgLItIDitbeN4rqjDgW01vv
sDaY6tTSS6ULZ/v1WReUkuryVj7cDoIlFqQ+gu6Osw2QXkGsZ/BuF2TxFSY92Rl/4cb0H80bDRQq
C0QU5DVAKXBnCYlZhPh294sZQPy4xPkNxM+43yIp9JfeQKMT/AxK90Cq/tcOGOBPhMJMdc+XAaXA
uQwW4sv6Dh+XJMoZLAPSSRuYRNkz2g5XLZW6+XneEiKgxJM0sdmFnvNhKy2JqGpCRiNo1ee0VL8J
bzsEuSq8r6PBoHrybmaxytH8yYSXezZGoCgB7GxHqskTmRh7aYkMStS51DFna9OrKciCSqpyc2E+
ElpYPeOhrld+DY0GziiSiYFDSWD34d6nXS2myPnd296+XRazoaI0HykMTWnLL0d75B+TsN3fSwKj
mEzSFs7plBM3ajlU8I31A8e5yMJzFuHa+xOTl9GoZaqskgv1OkWXhthmMckgdoPYruX6DTqMjxYr
LENVBZUZwMqztRbnB37hBgOgoZTVObG1eNsG+XSbBAn94tY3Y7CA9tF6Iu8lHi5oifh01mRc7qtQ
g7JGbQW8JurtG4s7AUNx8oC9jx/oBzF2iF1h6dObvBb7g7ZyJkYs9w6HOIYZqCtIxboLhliRnjn7
t48MThvf0ZCIc7Q4XAgCh0P0P8NBfPPRAwg+bLAkBQmsJkm8hhd1HeiDJNGIHBV99+2fFKNLgctM
X6Wq1eztjDYGnA8/8+ldJCnju29yOCZrXwC7iEODHF9xg5H+UcuR9bohO9lFVPBZV6kPWVq/s/kQ
XpGq3UH5Y+6lUhj/Oxr3XuxGtlmqFBz6Uc9hB9LouVYOGCthI6j2oXmqFEt3UgGgMtbgf2JXSpJD
9vCZOfhRciGDsVPJeaKyKcRebtQV0JqAV/waqLMH+AzggDAvW2g/jg81bIrUZO3ffclb3DXGpWzq
ZSjd0cRu6p9h15ac3+8HFYC6MtPWxEtObGFWtEHvBJM5gh2LK28CptZdMmFiBn9P41HW3jHVWBb2
p8KDWcOQWUn27RoQjIw3LaHMG32J6ST7AzwCbM+Kly0Ei2dSbjYOYfyIMa8bycPsZyuv2rbkPm4M
sEXdSLkpL6EC5r8Oe2QMm6lr62ETbLKGG/J5z5dDQvtd2rmxoLvv93waPcz+4i2HDNchfZKW2tkJ
T6x21LvheRNuIEI+qDS29/ylL5BlwSPKt8xdCLq5oT/xcWd8MUmz4+KDB39/Cn5yOdxIu2btkFic
jOTnuBVLHnP590y1zGEXliiYiW+Mony2TJdYdwEVuRhvUyz2WEw9nySXlZzKfe7JLp8rSMKjTGyz
CfFwL8firsd4oOpLrWdF5qGSZXI0KLQ3zQFHkQO/l/q5dAt/9YG9u8HV/J3tO3gPgoecee625MQb
/E4KBMtwq6CLJw/pcjP+HR46CcWzrlQyA7ho5LfrjslDZAza+RaCy/WfNw9B4Lx5nGaCdsLOjNJG
R08TEzVXqtxCqnBQ88cmvkCHVNoqon42bAqD67a24VEe+lo+NGdWuHqxSZ1A55d5AvaoB5A20ELX
5nnJgCkVwuy4Br2O/ub3PNOGAGJUj04v60bQqDy/UUmljAXwfDyIyxiTl8WuNlGqNb947kSHA97U
TPFR+LgXmyIwaQwsYWPf9vBzKtcyHs0udSr5avPlcP59TfWEzTdBRv/qkPBNJiorqOEQC5H6dlVs
q128nAAm3HGCYypaH5AZFVBuuIkgrr51EXB3BRib3gGUIPynQOo/+wdV/9/szWxF5KKaStN5zuUA
l0LSErPDXsr2QytMsv8cN0LFzD/+Pl+dWsPjam6wya2829owCS4bqa9fXrGl/ACRCmNi9v2T2WP2
qzbKtrfAsnbUvpao49KzGpi9l+tfsAT77+or0Cy7AxEn1emr4betT39m9ReoDz5dfQVRsgZtvLDF
xuQqtDCCf81wWJhRgEMerQDXlcAW14yQK9yhmZyEBjSgoB4M2YYi3AN7zm2EZEQF3oAQ6Sd+F1Ul
ml7N/pGdt82Ge8WTSRfasS+u1jxgikfdu8wqlgWBFskFm0We6NwWzSuqfyV2NjwGVFSG/K4zseG4
fZhZ4j0d9R5ObFXw0wOAKa/SPyZfhO5PwC2pjtWi6zsOibEyl3RNPfMReuN882UNPjRm77QE4ril
cMOMELFn3PMx3coD1+5ZBaa/rvFilk7Py5CPxdvjdGCwZ0M65XDYSRzjKu2MD09Qlrdi6Zb7QtIV
pAGzLG0ian+G2jVz+JoIhOWCJDobibL3buJ+6HGpQ7LSCX9xrsmiPLInDWKfLH0ZPvBcxOt0+hQr
IbGTABd1vSxgBH3P7rl376huEzGzGGsIZr6DPosWy/we2vnf/sRckfjFf/7FVvGqw/nihNMg5gr0
EeZrqhkWANsXttyTDiLFPRmoypmx2ehjbP/3deycIcn6YOV5/r5rPXQwKtUJGKhhfavz6BbMLrjN
z7w0mbxdOVesmttW7hb1Pfgu8nM0XOPw/bh+T5xOERmwws/cu2FcFpzq5HI3fL8WsbjQ50paHwxV
WNwAQHsyD98A4u8O7fFkXoQqYDKAiYfIJ5uH0tXbruilyadaHtzFBrJardhKvtLjIYfovZIlNc9+
T2JdHhd1O9PUTXvdgjHFuSHCGAVurhC3O47u/K0fck8FdxEedODaAq/w8y86qNJAhfrpFdvhYhWv
f/7c/RHuvajrI4lHszyL3irwiwnC7Cx4nWo2tMc/Kp/XmQWMW2EnyGBahVXbxKZd26qIh9GFJIZj
2lsbvBLqJ1FnKFmRn5QxA4BuOdx5ig1mEVSfr1m1uy/fLtW9Bd6f7RzETELfAYjAaM+k7RMCQSDA
lQrCDj2GHTtpJuzDnbbRU46ObnoR3BDiBrc+gnHV/1RLOqCRpB3Os61CH3sdIs2S29w1yr0tlOFD
4s99P5TAing4KsUmtLa8IqzTbKF8d7UVfUWfqhSIkHZB4WovFQ3pmIYVe+GNuuMHhUNrXnfYZmx7
/FttI1z5HutGzmxp0LXYLT61A8VRQh0v/VFkxVLhpQUqtAC0xPp+Hyt40ZXur0ry0yAmffKVDJX8
emV4nnmQ1dXGgGW/P3Gvri9F1bKDREIXsqPmfAORgGc3BmU42+kF0lcCvsHFSK8iaZICYdZ6s2j+
mT7tTWsIpyvkOXPnglX2ynW7I+LyB/wniZ2NbYv2KfvQ8aHQejYKfV9ujVlmsGvoUGBp+hv97zS9
vj7nF1vbIYRGdbyFcvNk5ORRpJnuj2kj/nW3pygMVJ+DP2dzOhJEtGbLNobovLqZ2UxeONorPyPT
p1plyoSyHa6hUUvl4I4IosQt6mHLsUMkrVmq8hPHe02hZG2zXaEDv7a0Em3JmHO0XpwmuvxhEYMN
wp1wQqsUG+Z5KdXDTHq5ykURAbOSHH5KoD/urwXy21VSTFW74yn6gpGxdycIPLKy7T3PpscuHjR3
yWUkQ/1aPYVonUuv0Wzven7aE3dCANN0kE2fBWNgIWRlpBye6dU2FpA2QAFUuHIyQeXvippZbP2L
4ysWUaqM2XXfUrmj2adjklb97Qy1dlAM4T/vVhPweiNBhKMnQxAfxPl0RCGcCFYUAZiOs8GZFTey
gEsPBlHhOllSYZh2dshsJ//4D+H60UFBXB1e5rC73Z3ty0XTn24m0lAZT4akT2Jza/TplSvJ1P30
AeflMvDhCUqyhOxdRgXzQ+KgtyI1YAvJHzKUnZgAuhRUMj1Wpj3/ISDVasmUBZxa4DE5jkRyywbM
it9Zjr7rSzTVNUJHk9v6FZMLIYSrQ4FS7YMYslydd23IoPmArWjnZoN+cKgCAKiIKTS7eK100ljL
b+74ALQTJ4TSy8XBUgMt44hKwKir5UeslDbsjLbIpKywsjxgypyvhE8iWNuAMJ1WVvMyW9Weauip
E4yaD6VSJ5h16pUmmmQsCQlf44g3nx1PVnw56ttaBdlwlV+S+zBBu80XjSfd5LitoeUSeNIgc+Ki
GD6A41OdkLSHR9F+D+3wFbR7l4CmsvuvW47EOj241YqSD9MRgbZWq5+DrtPH5r2jYxWun5YFo1KF
7ZEt20s3kNvcNJJkMHzLhqy6O4dSvJR7O40tXXcbxS9Fo3hVEh3QnDBPlGjSuP10KZJrytGDz2RP
hLwqUl37BLKqWuSou0mJR11inwIJsvOkMh//ODrplB5RjUONzCSq72PNKcFm05eA0RxAo5kIVIrg
mt/OUBV80O+vNwIa0RgooJj9k+DJuZT30zPIuqTjYrk6bhG+fpCx2Dw6XCh+yXXsErPx1cBGLZSE
pEkm29dGunL2Xr/cKziWKYgtSxKLJ6mboUwf0Y8PRcT2jctipR0lZxK3i/dw5r559lUBCjCG0EdG
Bs4gNYqhNlX90010MNnfUSMdjhtfoNO7dk4hdx7+IHxW2hKCmWqYBUAHVjKaN9nkWqiG/AyX72nv
4cFMunsz+ytHvpfX6sEZkvyr27qCnJTKLH5EkhVVLgPkPHe0hkAGMPQJBovGZlA46xsVvS2cX7+P
X8t6H15NNrzOlMFeuD/UyGMMtjsmmACjCI5lhNIM0kwrwMhJ9YNldVMC1u4O/kZhAbk2bvn99sWM
+5HcKyjiv84Y0mIJuNFtt95vpb7KNvNPy2IMFCzWd18qRum9bR3+inERLaOjecc7a5KK3xC4Ue8H
mCZyAs7R1IBOn4D+jtstQrkd6QyTYzT/5QDmlzdDrJtZV8zsi64DcSK2q7ynRa7Gc81hcHQsbVmF
s4s87d3zaOxpxV/Dwhe7HtQfkEvauF2iOtH3q9/9+3yulpQva53V+/YyOiAQH2F1ARLnGPy6KlZl
aY0Jo5wmYrlaFtvzviEBk2IWWzw4ZahO9KzH4XhZI0Ly3xOa4NkdzsgafZO/NCVhxc1bbQA1Qrfr
iIpqIadLg6bIT5E/V8+LTwLKERBKehGn5cup9ndU0b5G1w1hqlTXb+XwddByEAp2oK2g4IzzenXt
t/nAoq/S/X69/9HFjpf9HNhROxKF86w4rlzqnLmpxOfqJcfe43RgP1rgrJX2NHOU4ivJzXGGy+6S
ueuuTWSxY1UB4djmkff4Xna2I58OOlFgZ93BFNACNScwNuDm5sxH0WLoQ6i+hGIn9fFKi41Ili0b
8H4mAc5KIiB+7xf+T9YP/pYuq6e3n/qLnIQDHqVlnKjCtMeQQ70w0zro3vvL4MWEoxJ2uY/iIrTN
Nyxb7J/RUqY3eM0f7JpyESRfb4HE2LzDR2VYDkW72W0LHhcdDoPK5EpJ2VfpD6kP8EeGi+Rg4/xb
+vHuCB29vKNK3ZHShT3CjT+O9KvUrPyPuQhB6trcnQBnT7B7PLGBV08VNHq2H2RqUpzy8Q1qwyF+
+FQ/xkOyXFmCW6z7QWfCmsZuDUZZXlChZVZ8uVe0S1RyHXTLhpwRVK5K0Q8E33gwiwXsjwyJnX+F
AYLzh+a18FnE81gTZmUexlDvVlbG+xAP3bg9Bpo1xa+6IT3YoaGVTNCea1hKT0DrQDH3wykBu4Ez
d7/R78btABBKNkmNWkJ+AIBlhBZMh4HTBLthIm8vBkeDrxOgHCJdTralOvwN0PtADvYM1s26
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity vga_dvi_tx is
port(
  I_rst_n :  in std_logic;
  I_serial_clk :  in std_logic;
  I_rgb_clk :  in std_logic;
  I_rgb_vs :  in std_logic;
  I_rgb_hs :  in std_logic;
  I_rgb_de :  in std_logic;
  I_rgb_r :  in std_logic_vector(7 downto 0);
  I_rgb_g :  in std_logic_vector(7 downto 0);
  I_rgb_b :  in std_logic_vector(7 downto 0);
  O_tmds_clk_p :  out std_logic;
  O_tmds_clk_n :  out std_logic;
  O_tmds_data_p :  out std_logic_vector(2 downto 0);
  O_tmds_data_n :  out std_logic_vector(2 downto 0));
end vga_dvi_tx;
architecture beh of vga_dvi_tx is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
component \~rgb2dvi.vga_dvi_tx\
port(
  I_rgb_clk: in std_logic;
  I_serial_clk: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  I_rst_n: in std_logic;
  I_rgb_de: in std_logic;
  I_rgb_vs: in std_logic;
  I_rgb_hs: in std_logic;
  I_rgb_r : in std_logic_vector(7 downto 0);
  I_rgb_g : in std_logic_vector(7 downto 0);
  I_rgb_b : in std_logic_vector(7 downto 0);
  O_tmds_clk_p: out std_logic;
  O_tmds_clk_n: out std_logic;
  O_tmds_data_p : out std_logic_vector(2 downto 0);
  O_tmds_data_n : out std_logic_vector(2 downto 0));
end component;
begin
GND_s3: GND
port map (
  G => GND_0);
VCC_s3: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
rgb2dvi_inst: \~rgb2dvi.vga_dvi_tx\
port map(
  I_rgb_clk => I_rgb_clk,
  I_serial_clk => I_serial_clk,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  I_rst_n => I_rst_n,
  I_rgb_de => I_rgb_de,
  I_rgb_vs => I_rgb_vs,
  I_rgb_hs => I_rgb_hs,
  I_rgb_r(7 downto 0) => I_rgb_r(7 downto 0),
  I_rgb_g(7 downto 0) => I_rgb_g(7 downto 0),
  I_rgb_b(7 downto 0) => I_rgb_b(7 downto 0),
  O_tmds_clk_p => O_tmds_clk_p,
  O_tmds_clk_n => O_tmds_clk_n,
  O_tmds_data_p(2 downto 0) => O_tmds_data_p(2 downto 0),
  O_tmds_data_n(2 downto 0) => O_tmds_data_n(2 downto 0));
end beh;
