--Copyright (C)2014-2024 Gowin Semiconductor Corporation.
--All rights reserved.
--File Title: IP file
--Tool Version: V1.9.10 (64-bit)
--Part Number: GW2A-LV18PG256C8/I7
--Device: GW2A-18
--Device Version: C
--Created Time: Mon Jul 22 14:34:06 2024

library IEEE;
use IEEE.std_logic_1164.all;

entity VGA_FONT_pROM is
    port (
        dout: out std_logic_vector(7 downto 0);
        clk: in std_logic;
        oce: in std_logic;
        ce: in std_logic;
        reset: in std_logic;
        ad: in std_logic_vector(11 downto 0)
    );
end VGA_FONT_pROM;

architecture Behavioral of VGA_FONT_pROM is

    signal prom_inst_0_dout_w: std_logic_vector(27 downto 0);
    signal prom_inst_1_dout_w: std_logic_vector(27 downto 0);
    signal gw_gnd: std_logic;
    signal prom_inst_0_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_0_DO_o: std_logic_vector(31 downto 0);
    signal prom_inst_1_AD_i: std_logic_vector(13 downto 0);
    signal prom_inst_1_DO_o: std_logic_vector(31 downto 0);

    --component declaration
    component pROM
        generic (
            READ_MODE: in bit :='0';
            BIT_WIDTH: in integer := 1;
            RESET_MODE: in string := "SYNC";
            INIT_RAM_00: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_01: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_02: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_03: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_04: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_05: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_06: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_07: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_08: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_09: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_0F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_10: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_11: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_12: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_13: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_14: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_15: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_16: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_17: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_18: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_19: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_1F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_20: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_21: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_22: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_23: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_24: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_25: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_26: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_27: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_28: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_29: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_2F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_30: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_31: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_32: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_33: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_34: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_35: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_36: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_37: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_38: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_39: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3A: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3B: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3C: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3D: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3E: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000";
            INIT_RAM_3F: in bit_vector := X"0000000000000000000000000000000000000000000000000000000000000000"
        );
        port (
            DO: out std_logic_vector(31 downto 0);
            CLK: in std_logic;
            OCE: in std_logic;
            CE: in std_logic;
            RESET: in std_logic;
            AD: in std_logic_vector(13 downto 0)
        );
    end component;

begin
    gw_gnd <= '0';

    prom_inst_0_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(3 downto 0) <= prom_inst_0_DO_o(3 downto 0) ;
    prom_inst_0_dout_w(27 downto 0) <= prom_inst_0_DO_o(31 downto 4) ;
    prom_inst_1_AD_i <= ad(11 downto 0) & gw_gnd & gw_gnd;
    dout(7 downto 4) <= prom_inst_1_DO_o(3 downto 0) ;
    prom_inst_1_dout_w(27 downto 0) <= prom_inst_1_DO_o(31 downto 4) ;

    prom_inst_0: pROM
        generic map (
            READ_MODE   => '0',
            BIT_WIDTH   => 4,
            RESET_MODE  => "SYNC",
            INIT_RAM_00 => X"000008CEEEEC00000000EFF73FFBFE000000E119D1151E000000000000000000",
            INIT_RAM_01 => X"0000008CC80000000000C88EFFEC80000000C88777CC80000000008CEC800000",
            INIT_RAM_02 => X"00008CCCC82AEE00FFFFF39DD93FFFFF00000C6226C00000FFFFFF7337FFFFFF",
            INIT_RAM_03 => X"000088BC7CB8800000006773333F3F0000000000000F3F00000088E8C6666C00",
            INIT_RAM_04 => X"0000660666666600000008CE888EC800000026EEEEEEE620000000008E800000",
            INIT_RAM_05 => X"0000E8CE888EC8000000EEEE00000000000C6C8C66C806C00000BBBBBBBBBF00",
            INIT_RAM_06 => X"00000000E00000000000008CEC80000000008CE88888880000008888888EC800",
            INIT_RAM_07 => X"00000088CCEE000000000EECC88000000000008CEC800000000000E000000000",
            INIT_RAM_08 => X"0000CCECCCECC00000000000000466600000880888CCC8000000000000000000",
            INIT_RAM_09 => X"000000000000000000006CCCC68CC800000066008C6200000088C6666C026C88",
            INIT_RAM_0A => X"00000088E88000000000006CFC600000000008CCCCCC80000000C80000008C00",
            INIT_RAM_0B => X"000000008C620000000088000000000000000000E00000000000888000000000",
            INIT_RAM_0C => X"0000C6666C666C000000E60008C66C000000E8888888880000008C666666C800",
            INIT_RAM_0D => X"000000008C666E000000C6666C0008000000C6666C000E000000ECCCECCCCC00",
            INIT_RAM_0E => X"0000088000880000000008800088000000008C666E666C000000C6666C666C00",
            INIT_RAM_0F => X"0000880888C66C000000008C6C8000000000000E00E0000000006C80008C6000",
            INIT_RAM_10 => X"0000C62000026C000000C6666C666C0000006666E66C80000000C0CEEE66C000",
            INIT_RAM_11 => X"0000A666E0026C000000000088826E000000E62088826E0000008C666666C800",
            INIT_RAM_12 => X"0000666C88C6660000008CCCCCCCCE000000C88888888C00000066666E666600",
            INIT_RAM_13 => X"0000C66666666C0000006666EEE666000000666666EEE6000000E62000000000",
            INIT_RAM_14 => X"0000C666C8066C0000006666CC666C0000ECCE6666666C00000000000C666C00",
            INIT_RAM_15 => X"0000CEE666666600000008C6666666000000C666666666000000C888888AEE00",
            INIT_RAM_16 => X"0000C00000000C000000E62008C66E000000C8888C666600000066CC88CC6600",
            INIT_RAM_17 => X"00F00000000000000000000000006C800000CCCCCCCCCC00000026EC80000000",
            INIT_RAM_18 => X"0000C60006C000000000C6666C80000000006CCCCC8000000000000000000800",
            INIT_RAM_19 => X"08CCCCCCCC600000000000000004C8000000C600E6C0000000006CCCCCCCCC00",
            INIT_RAM_1A => X"000066C88C6000000C66666666E066000000C888888088000000666666C00000",
            INIT_RAM_1B => X"0000C66666C000000000666666C00000000066666EC000000000C88888888800",
            INIT_RAM_1C => X"0000C6C806C000000000000066C000000ECCCCCCCC6000000000C66666C00000",
            INIT_RAM_1D => X"0000CE666660000000008C666660000000006CCCCCC000000000C60000C00000",
            INIT_RAM_1E => X"0000E88880888E000000E6008CE0000008C6E6666660000000006C888C600000",
            INIT_RAM_1F => X"00000E666C800000000000000000C600000008888E8880000000888880888800",
            INIT_RAM_20 => X"00006CCCCC80C8000000C600E6C008C000006CCCCCC00C0000C6CC6200026C00",
            INIT_RAM_21 => X"000C6CC6006C000000006CCCCC808C8000006CCCCC80800000006CCCCC800C00",
            INIT_RAM_22 => X"0000C888888006000000C600E6C080000000C600E6C006000000C600E6C0C800",
            INIT_RAM_23 => X"0000666E66C808C80000666E66C800600000C888888080000000C88888806C80",
            INIT_RAM_24 => X"0000C66666C0C8000000ECCCCECCCE000000E88E66C000000000E600C06E0008",
            INIT_RAM_25 => X"00006CCCCCC0800000006CCCCCC0C8000000C66666C080000000C66666C00600",
            INIT_RAM_26 => X"000088C60006C8800000C666666660600000C6666666C06008C6E66666600600",
            INIT_RAM_27 => X"000888888E888BE000006CCCEC48CC800000888E8E8C66000000C60000004C80",
            INIT_RAM_28 => X"00006CCCCCC000800000C66666C000800000C888888008C000006CCCCC800080",
            INIT_RAM_29 => X"000000000C08CC80000000000E0ECCC00000666EEE6660C60000666666C0C600",
            INIT_RAM_2A => X"00E8C6C008C62000000006666E000000000000000E0000000000C66000000000",
            INIT_RAM_2B => X"0000008C6C8000000000006C8C60000000008CCC888088000066EEE608C62000",
            INIT_RAM_2C => X"88888888888888887D7D7D7D7D7D7D7DA5A5A5A5A5A5A5A54141414141414141",
            INIT_RAM_2D => X"66666666E0000000666666666666666688888888888888888888888888888888",
            INIT_RAM_2E => X"6666666666E00000666666666666666666666666666666668888888888800000",
            INIT_RAM_2F => X"8888888880000000000000008888888800000000E666666600000000E6666666",
            INIT_RAM_30 => X"88888888F888888888888888F000000000000000F888888800000000F8888888",
            INIT_RAM_31 => X"666666667666666688888888F8F8888888888888F888888800000000F0000000",
            INIT_RAM_32 => X"6666666670F0000000000000F07666666666666670F0000000000000F0766666",
            INIT_RAM_33 => X"00000000F0F88888666666667076666600000000F0F000006666666670766666",
            INIT_RAM_34 => X"00000000F666666666666666F000000088888888F0F0000000000000F6666666",
            INIT_RAM_35 => X"66666666F666666666666666F000000088888888F8F0000000000000F8F88888",
            INIT_RAM_36 => X"FFFFFFFFFFFFFFFF88888888F0000000000000008888888888888888F8F88888",
            INIT_RAM_37 => X"000000000FFFFFFFFFFFFFFFFFFFFFFF0000000000000000FFFFFFFFF0000000",
            INIT_RAM_38 => X"0000CCCCCCCE00000000000000066E000000C666C8CCC80000006C888C600000",
            INIT_RAM_39 => X"0000888888C60000000000C6666600000000088888E000000000E6008006E000",
            INIT_RAM_3A => X"0000C6666EC80E000000ECCCC666C80000008C66E66C80000000E8C666C8E000",
            INIT_RAM_3B => X"000066666666C0000000C0000C000C00000000E3BBE63000000000EBBBE00000",
            INIT_RAM_3C => X"0000E0C80008C0000000E008C6C800000000F0088E88000000000E00E00E0000",
            INIT_RAM_3D => X"000000C60C60000000000880E0880000000008888888888888888888888BBE00",
            INIT_RAM_3E => X"0000CCCCCCCCCCF000000008000000000000000880000000000000000008CC80",
            INIT_RAM_3F => X"000000000000000000000CCCCCCC00000000000008800800000000000CCCCC80"
        )
        port map (
            DO => prom_inst_0_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_0_AD_i
        );

    prom_inst_1: pROM
        generic map (
            READ_MODE   => '0',
            BIT_WIDTH   => 4,
            RESET_MODE  => "SYNC",
            INIT_RAM_00 => X"0000137FFFF6000000007FFECFFDF70000007889B88A87000000000000000000",
            INIT_RAM_01 => X"000000133100000000003117FF7310000000311EEE33100000000137F7310000",
            INIT_RAM_02 => X"00007CCCC7310100FFFFFC9BB9CFFFFF0000036446300000FFFFFFECCEFFFFFF",
            INIT_RAM_03 => X"000011D3E3D11000000CEE66666767000000EF73333333000000117136666300",
            INIT_RAM_04 => X"00006606666666000000013711173100000000013F31000000008CEFFFFFEC80",
            INIT_RAM_05 => X"00007137111731000000FFFF000000000007C036CC636C700000111117DDD700",
            INIT_RAM_06 => X"00000036F630000000000010F010000000001371111111000000111111173100",
            INIT_RAM_07 => X"0000013377FF000000000FF77331000000000026F6200000000000FCCC000000",
            INIT_RAM_08 => X"000066F666F66000000000000002666000001101113331000000000000000000",
            INIT_RAM_09 => X"000000000006333000007CCCD736630000008C6310CC000000117C8007CCC711",
            INIT_RAM_0A => X"000000117110000000000063F360000000003100000013000000013333331000",
            INIT_RAM_0B => X"00008C6310000000000011000000000000000000F00000000003111000000000",
            INIT_RAM_0C => X"00007C000300C7000000FCC63100C7000000711111173100000036CCDDCC6300",
            INIT_RAM_0D => X"000033331000CF0000007CCCCFCC630000007C000FCCCF0000001000FC631000",
            INIT_RAM_0E => X"000031100011000000000110001100000000700007CCC70000007CCCC7CCC700",
            INIT_RAM_0F => X"00001101110CC700000063100013600000000007007000000000001363100000",
            INIT_RAM_10 => X"000036CCCCCC63000000F66667666F000000CCCCFCC6310000007CDDDDCC7000",
            INIT_RAM_11 => X"000036CCDCCC63000000F66667666F000000F66667666F000000F66666666F00",
            INIT_RAM_12 => X"0000E66677666E0000007CCC0000010000003111111113000000CCCCCFCCCC00",
            INIT_RAM_13 => X"00007CCCCCCCC7000000CCCCCDFFEC000000CCCCCDFFEC000000F66666666F00",
            INIT_RAM_14 => X"00007CC0036CC7000000E66667666F0000007DDCCCCCC7000000F66667666F00",
            INIT_RAM_15 => X"00006EFDDDCCCC000000136CCCCCCC0000007CCCCCCCCC000000311111157700",
            INIT_RAM_16 => X"00003333333333000000FCC63108CF0000003111136666000000CC673376CC00",
            INIT_RAM_17 => X"00F0000000000000000000000000C63100003000000003000000000137EC8000",
            INIT_RAM_18 => X"00007CCCCC7000000000766666766E0000007CCC707000000000000000000133",
            INIT_RAM_19 => X"07C07CCCCC7000000000F6666F66630000007CCCFC70000000007CCCC6300100",
            INIT_RAM_1A => X"0000E66776666E00036600000000000000003111113011000000E66667666E00",
            INIT_RAM_1B => X"00007CCCCC7000000000666666D000000000CDDDDFE000000000311111111300",
            INIT_RAM_1C => X"00007C036C7000000000F66667D0000001007CCCCC7000000F66766666D00000",
            INIT_RAM_1D => X"00006FDDDCC00000000013666660000000007CCCCCC000000000133333F33100",
            INIT_RAM_1E => X"00000111171110000000FC631CF000000F007CCCCCC000000000C63336C00000",
            INIT_RAM_1F => X"00000FCCC6310000000000000000D70000007111101117000000111110111100",
            INIT_RAM_20 => X"00007CCC7070631000007CCCFC70310000007CCCCCC00C000070036CCCCC6300",
            INIT_RAM_21 => X"000300366663000000007CCC7070363000007CCC7070136000007CCC70700C00",
            INIT_RAM_22 => X"000031111130060000007CCCFC70136000007CCCFC700C0000007CCCFC706310",
            INIT_RAM_23 => X"0000CCCFCC6303630000CCCFCC6310C000003111113013600000311111306310",
            INIT_RAM_24 => X"00007CCCCC7063100000CCCCCFCC630000006DD737C000000000F666766F0631",
            INIT_RAM_25 => X"00007CCCCCC0136000007CCCCCC0C73000007CCCCC70136000007CCCCC700C00",
            INIT_RAM_26 => X"000011366666311000007CCCCCCCC0C000007CCCCCCC70C007007CCCCCC00C00",
            INIT_RAM_27 => X"007D1111171111000000CCCCDCCFCCF000001117171366000000FE6666F66630",
            INIT_RAM_28 => X"00007CCCCCC0631000007CCCCC706310000031111130310000007CCC70706310",
            INIT_RAM_29 => X"000000000703663000000000070366300000CCCCDFFEC0D70000666666D0D700",
            INIT_RAM_2A => X"003108D631CCCCC0000000000F00000000000CCCCF00000000007CCC63303300",
            INIT_RAM_2B => X"000000D636D0000000000036D63000000000133311101100000039C631CCCCC0",
            INIT_RAM_2C => X"11111111111111117D7D7D7D7D7D7D7DA5A5A5A5A5A5A5A54141414141414141",
            INIT_RAM_2D => X"33333333F000000033333333F333333311111111F1F1111111111111F1111111",
            INIT_RAM_2E => X"33333333F0F00000333333333333333333333333F0F3333311111111F1F00000",
            INIT_RAM_2F => X"11111111F000000000000000F1F1111100000000F333333300000000F0F33333",
            INIT_RAM_30 => X"111111111111111111111111F000000000000000F11111110000000011111111",
            INIT_RAM_31 => X"3333333333333333111111111111111111111111F111111100000000F0000000",
            INIT_RAM_32 => X"33333333F0F0000000000000F0F3333333333333333000000000000033333333",
            INIT_RAM_33 => X"00000000F0F1111133333333F0F3333300000000F0F000003333333333333333",
            INIT_RAM_34 => X"000000003333333333333333F000000011111111F0F0000000000000F3333333",
            INIT_RAM_35 => X"33333333F3333333333333333000000011111111111000000000000011111111",
            INIT_RAM_36 => X"FFFFFFFFFFFFFFFF111111111000000000000000F111111111111111F1F11111",
            INIT_RAM_37 => X"000000000FFFFFFF0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFF0000000",
            INIT_RAM_38 => X"00006666666F00000000CCCCCCCCCF000000CCCCCDCCC70000007DDDDD700000",
            INIT_RAM_39 => X"0000111111D70000000C66766666000000007DDDDD7000000000FC63136CF000",
            INIT_RAM_3A => X"00003666630131000000E6666CCC6300000036CCFCC630000000713666317000",
            INIT_RAM_3B => X"0000CCCCCCCC700000001366676631000000C67FDD7000000000007DDD700000",
            INIT_RAM_3C => X"000070013631000000007031000130000000F0011711000000000F00F00F0000",
            INIT_RAM_3D => X"000000D70D700000000001107011000000007DDD111111111111111111111000",
            INIT_RAM_3E => X"00001366E0000000000000010000000000000001100000000000000000036630",
            INIT_RAM_3F => X"00000000000000000000077777770000000000000FC63D7000000000066666D0"
        )
        port map (
            DO => prom_inst_1_DO_o,
            CLK => clk,
            OCE => oce,
            CE => ce,
            RESET => reset,
            AD => prom_inst_1_AD_i
        );

end Behavioral; --VGA_FONT_pROM
